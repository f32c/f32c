--
-- Copyright 2008, 2010 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
--

-- $Id: bram.vhd 116 2011-03-28 12:43:12Z marko $

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library xp2;
use xp2.components.all;


entity bram is
	generic(
		mem_type: string := "big"
	);
	port(
		clk: in std_logic;
		imem_addr: in std_logic_vector(31 downto 2);
		imem_data_out: out std_logic_vector(31 downto 0);
		imem_addr_strobe: in std_logic;
		imem_data_ready: out std_logic;
		dmem_addr: in std_logic_vector(31 downto 2);
		dmem_data_in: in std_logic_vector(31 downto 0);
		dmem_data_out: out std_logic_vector(31 downto 0);
		dmem_byte_we: in std_logic_vector(3 downto 0);
		dmem_addr_strobe: in std_logic;
		dmem_data_ready: out std_logic
	);
end bram;

architecture Behavioral of bram is
	signal dmem_wait_cycle, dmem_must_wait, dmem_we: std_logic;
	signal dmem_data_read, dmem_write_out: std_logic_vector(31 downto 0);
	signal dmem_bram_cs: std_logic;
begin
	
	imem_data_ready <= '1';
	dmem_data_out <= dmem_data_read; -- shut up compiler errors
	
	dmem_data_ready <= '1';
	dmem_write_out <= dmem_data_in;
	dmem_bram_cs <= dmem_addr_strobe;

	ram_0: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B=> "NORMAL", WRITEMODE_A => "NORMAL",
		GSR=> "DISABLED", RESETMODE=> "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A=> "NOREG",
		DATA_WIDTH_B=> 9, DATA_WIDTH_A=> 9,
		INITVAL_00 => "0x1FE00000070422104680000fb008210002110001104fc000110062502404000f9008000100114000",
		INITVAL_01 => "0x000070422310001000fd0080004221042800080010421000fc000150060002C0400008002fb00001",
		INITVAL_02 => "0x010ff010011F2ff00800006030062100008002fd0000104205000210140300008002fd000ff00600",
		INITVAL_03 => "0x00223000f3004f5080f7100420022b0044204A1104073042c00422100008084fa080210000200221",
		INITVAL_04 => "0x04280042230460010021046c00464010080020100D41d002240B61c006e018000010000000204Af1",
		INITVAL_05 => "0x0060006001042100426a01421020b7042210461c04024030d804008180211FEff0380404680046c0",
		INITVAL_06 => "0x1FE01010e204201002b30460005A280101803820048f8056ff0000100000000201A2240082b000f5",
		INITVAL_07 => "0x000730C625042210203c07034058180382004828068d000008002f71FE01000f7014300AE020020b",
		INITVAL_08 => "0x1FE001C2100900400030010180382004828042211FE10016011F02600200002fb002000580e00207",
		INITVAL_09 => "0x0380d04804048261901018800008011F44008421000fb00208080421F0010420e04218038141C021",
		INITVAL_0A => "0x04202070210004e008300100c1E0ac000000002001014030010400802818038ef05423008000A8c4",
		INITVAL_0B => "0x018001F82a04604000130080c00408018001DE01000fc0542300804018001F82a046040080c01003",
		INITVAL_0C => "0x000fc1102300804018020100000801006ff00000000101A001030c3000ac002fc054230080002604",
		INITVAL_0D => "0x0002100000006001C0000087b00C61006090060004214000c40002e05614042001F888046040080c",
		INITVAL_0E => "0x0200800808018bb008c41AA1405604000dd002001F888046040080c000fc11023008040180804A24",
		INITVAL_0F => "0x042f80428000000160251E0b004233038200482c06034050c800000042c007E2318001182dd00006",
		INITVAL_10 => "0x0200407008038200482805830068081F407018240420002A210427c046c008001106000282604021",
		INITVAL_11 => "0x042211A048040240501805821042140001c042d010028160fa04A0f000b000013042080421004248",
		INITVAL_12 => "0x028180382004828058000AAe8042081D8b8168ec1700104201010b403004158021440311A0104208",
		INITVAL_13 => "0x046210900004208042210421408623042481800700021070140283c1F41404C14040210A0e406008",
		INITVAL_14 => "0x000440420d002210D4600780400608042c0000231582618623026000002104240042080422105043",
		INITVAL_15 => "0x002ec042b40062113E88042021D8b4058a71B821018ec16864142000602102818038200482805864",
		INITVAL_16 => "0x1D8210587d04621180f4028211D801042ec042c4142041D8b4000f1058911E821168ec004961E821",
		INITVAL_17 => "0x1680e1D801168b41D82101Cc3000870C8a101Cec080010280e1D88304214046a118014008ec00204",
		INITVAL_18 => "0x17808006011780f04826020c4190211F61404C14040210A01c030d0028e00000000023142c01FE14",
		INITVAL_19 => "0x00061040750406f0CA6e0EC200CC730E66f040201882e040140301c04220178c405C14040140301c",
		INITVAL_1A => "0x0DC630D66f088740A6720B46908E000DE4b0CA5a0DE690DE530EC560CA750DC700406f0CA6c0EA20",
		INITVAL_1B => "0x0A8370900008040060da05014000ec1B0c41A8941808007E10000000DC670DE790C8200DC7a0DE20",
		INITVAL_1C => "0x000000000000000000000000000000000a000498008900108800480008780107d0D89a0C81f0B8c9",
		INITVAL_1D => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DIA0 => dmem_write_out(0), DIA1 => dmem_write_out(1),
		DIA2 => dmem_write_out(2), DIA3 => dmem_write_out(3),
		DIA4 => dmem_write_out(4), DIA5 => dmem_write_out(5),
		DIA6 => dmem_write_out(6), DIA7 => dmem_write_out(7),
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(0), DOA1 => dmem_data_read(1),
		DOA2 => dmem_data_read(2), DOA3 => dmem_data_read(3),
		DOA4 => dmem_data_read(4), DOA5 => dmem_data_read(5),
		DOA6 => dmem_data_read(6), DOA7 => dmem_data_read(7),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => dmem_addr(2), ADA4 => dmem_addr(3),
		ADA5 => dmem_addr(4), ADA6 => dmem_addr(5),
		ADA7 => dmem_addr(6), ADA8 => dmem_addr(7),
		ADA9 => dmem_addr(8), ADA10 => dmem_addr(9),
		ADA11 => dmem_addr(10), ADA12 => dmem_addr(11),
		ADA13 => dmem_addr(12),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_byte_we(0),
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(0), DOB1 => imem_data_out(1),
		DOB2 => imem_data_out(2), DOB3 => imem_data_out(3),
		DOB4 => imem_data_out(4), DOB5 => imem_data_out(5),
		DOB6 => imem_data_out(6), DOB7 => imem_data_out(7),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => imem_addr(2), ADB4 => imem_addr(3),
		ADB5 => imem_addr(4), ADB6 => imem_addr(5),
		ADB7 => imem_addr(6), ADB8 => imem_addr(7),
		ADB9 => imem_addr(8), ADB10 => imem_addr(9),
		ADB11 => imem_addr(10), ADB12 => imem_addr(11),
		ADB13 => imem_addr(12),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_1: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B=> "NORMAL", WRITEMODE_A => "NORMAL",
		GSR=> "DISABLED", RESETMODE=> "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A=> "NOREG",
		DATA_WIDTH_B=> 9, DATA_WIDTH_A=> 9,
		INITVAL_00 => "0x1FE00000000402806048000ff000180001808000090ff000000001000000000ff000e00060011A00",
		INITVAL_01 => "0x000000403009000000ff0000002018070400003c09010024ff00000000000000000000000ff00000",
		INITVAL_02 => "0x000ff000001FE0000000034000001000000000ff0000002000000180000000000000ff000ff05C2e",
		INITVAL_03 => "0x00020000ff000ff020ff09E40000500001805000000000202f0701800000050ff040100000000010",
		INITVAL_04 => "0x0202803028040310702005021050310522000000000f3000d900E00000ff100000000000000050ff",
		INITVAL_05 => "0x03C1e0000004000060000008800000110800000000000000ff00000100101FE7f000000201003020",
		INITVAL_06 => "0x1FE0000000030000000004000000000000000000000ff030ff0000000000000000000000020000ff",
		INITVAL_07 => "0x0000000000110800000000000000000000000000000ff00000000ff1FE00042ff000000001700000",
		INITVAL_08 => "0x000001FE0000000000000000000000000000208800000000001FE1800000000ff000000000000000",
		INITVAL_09 => "0x0000003000040201008010000000001FE1003080000ff0000002018048001000002000000001FE88",
		INITVAL_0A => "0x07000000280400000000000001FE80000000000000000000000000000000000ff020100000000280",
		INITVAL_0B => "0x000001FE1002000110000000000000000001FE00000ff0301800000000001FE18030000000000000",
		INITVAL_0C => "0x000ff0261000000000000000000000000f90040400C00100001006800080000ff020100008800000",
		INITVAL_0D => "0x00C0000C0003C1e1FE0000000000000540003C1e04080000800000002000070001FE130200000000",
		INITVAL_0E => "0x0000000000000ff000801FE8002000000ff000001FE130200000000000ff02610000000000006030",
		INITVAL_0F => "0x120801209002200100100008013000000000000000000000ff000000E00100070002001FEff00000",
		INITVAL_10 => "0x0000000000000000000000000000001FE00000100500000080110801101011200020000000000020",
		INITVAL_11 => "0x04030100000000000000000201000000000020ff0208010001020000328000002060000400004000",
		INITVAL_12 => "0x00000000000000000000000030020000280100011000004000000800000000000000000000005000",
		INITVAL_13 => "0x05020000001300004030050000502804000120000001000000100801FE0000000000200008000000",
		INITVAL_14 => "0x0000002000000300003400400000000500c000200002002E20102000009010080040000503000028",
		INITVAL_15 => "0x0000105080000801FE130020000280000ff00A010000110000004000000100000000000000000000",
		INITVAL_16 => "0x00220000ff0400104001100280020005001040090040000280000ff000ff0020110001000ff00201",
		INITVAL_17 => "0x10000002001008000220000280000000002000010500010000002280408004002040800000100000",
		INITVAL_18 => "0x1000000000100000301810080100201FE0000000000200000000080000ff00000000200041000280",
		INITVAL_19 => "0x000660E663040720DA690C2500DE650D66d0826b1000200000000000400310080004800000000000",
		INITVAL_1A => "0x0DE72000760EA000E0000C2630DE000EC610C4610C8200DC6c0C275000630CA6c040720DA690C850",
		INITVAL_1B => "0x01A0001A0001Aff01Afe01A0d01A0c0180c00000000000000000000000720EE65000200DE650007a",
		INITVAL_1C => "0x0000000000000000000000000000000000d0000d0000d0000d0000d0000d0000201A0101A0101A00",
		INITVAL_1D => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DIA0 => dmem_write_out(8), DIA1 => dmem_write_out(9),
		DIA2 => dmem_write_out(10), DIA3 => dmem_write_out(11),
		DIA4 => dmem_write_out(12), DIA5 => dmem_write_out(13),
		DIA6 => dmem_write_out(14), DIA7 => dmem_write_out(15),
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(8), DOA1 => dmem_data_read(9),
		DOA2 => dmem_data_read(10), DOA3 => dmem_data_read(11),
		DOA4 => dmem_data_read(12), DOA5 => dmem_data_read(13),
		DOA6 => dmem_data_read(14), DOA7 => dmem_data_read(15),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => dmem_addr(2), ADA4 => dmem_addr(3),
		ADA5 => dmem_addr(4), ADA6 => dmem_addr(5),
		ADA7 => dmem_addr(6), ADA8 => dmem_addr(7),
		ADA9 => dmem_addr(8), ADA10 => dmem_addr(9),
		ADA11 => dmem_addr(10), ADA12 => dmem_addr(11),
		ADA13 => dmem_addr(12),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_byte_we(1),
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(8), DOB1 => imem_data_out(9),
		DOB2 => imem_data_out(10), DOB3 => imem_data_out(11),
		DOB4 => imem_data_out(12), DOB5 => imem_data_out(13),
		DOB6 => imem_data_out(14), DOB7 => imem_data_out(15),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => imem_addr(2), ADB4 => imem_addr(3),
		ADB5 => imem_addr(4), ADB6 => imem_addr(5),
		ADB7 => imem_addr(6), ADB8 => imem_addr(7),
		ADB9 => imem_addr(8), ADB10 => imem_addr(9),
		ADB11 => imem_addr(10), ADB12 => imem_addr(11),
		ADB13 => imem_addr(12),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_2: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B=> "NORMAL", WRITEMODE_A => "NORMAL",
		GSR=> "DISABLED", RESETMODE=> "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A=> "NOREG",
		DATA_WIDTH_B=> 9, DATA_WIDTH_A=> 9,
		INITVAL_00 => "0x18C82000c0104a2192090CE48084a20CE820102800Cc600040084a4080c2000000F41b0001d1381c",
		INITVAL_01 => "0x000c0112c8012290004308447100681C4091060200C4500Ac60004010400080c2000e014Ac014484",
		INITVAL_02 => "0x100421C0421406510883006a008A00000e00846010684000601060008082000e0108c010Ac600A05",
		INITVAL_03 => "0x08485000400D4a000440012051CE850D203050eb0160000005000a0000e000A80008440006014600",
		INITVAL_04 => "0x14405106e51880400Ac4144031480300402146a6000a500A84008bf100bd108001C0c4000c0050eb",
		INITVAL_05 => "0x006030C622080a30800000A4016400000a0100b1164bf160bd17Ae0104430C60317E410C40210603",
		INITVAL_06 => "0x14E6301000000a516000008a2004bd1C0b0162b217E60022310481000604046b2000bf1001104680",
		INITVAL_07 => "0x004140261200080144a714Ca517Eb0162b2166b4144bd000e014A6814C63008400844608E0414A68",
		INITVAL_08 => "0x00000080a200042088bd1C0b0162b2166b404023000a20A8630A65202002020520620217E4002052",
		INITVAL_09 => "0x17E600C4801064410483108620E2640800200602000800C840004030C60300080100b117Eb017A22",
		INITVAL_0A => "0x00008012000840216040162b217A8200000000bd1C0b01620217Ae0160b117E400A0510C40000082",
		INITVAL_0B => "0x0C40008043088620C6030C862004620040014Ca5000600C4640C6640CE000C0620C8630C8680D206",
		INITVAL_0C => "0x00040084430C4630C4020C402010090140b032180181111Ead1200d0DA8200440086440C46300664",
		INITVAL_0D => "0x1A44c08462006030C600080620806200Aa0006050008e1CA86000401DEef1C00008042086620C662",
		INITVAL_0E => "0x17Ae0160b116411020860808e1DEe7000881080008042086620C66900040084430C4630D46308Ccb",
		INITVAL_0F => "0x084820840400862104a20848214080160b1164b416Abf166bd000001A4001A4d2000521A45900058",
		INITVAL_10 => "0x14A3517Ae0160b1164b3168b517E3102810080620A022028000468304402004420046200C0000A40",
		INITVAL_11 => "0x0804012200166b416Ab117E40100b00A4b20C4bd00883104000C44200A820000008000140a514000",
		INITVAL_12 => "0x160b1164b3168b517E0008004000050008410400106430804200A820040200402004020040204000",
		INITVAL_13 => "0x10460000730E4001404004Aa500A8214000024520AA700A01412493024060001000A000649017Ae0",
		INITVAL_14 => "0x0C4020004008400000a500A6400C000808400882000440088210A04084520A0820C00004A4014A05",
		INITVAL_15 => "0x02000000840220008004000050008417E400080000A00108040006217A00160b1164b3168b517E04",
		INITVAL_16 => "0x0000017E4000800008101080000004000000000400005000840001117E40008001080000A4000800",
		INITVAL_17 => "0x108a50000410A820000014A02000000080014A0000A0410Aa50000500085008000088400A0000805",
		INITVAL_18 => "0x1086010684108600C8431088310400022060001000A00022bf16290160bd00000000820000210882",
		INITVAL_19 => "0x0006f0CA6e040000C2200E46f0E46d0D2610EA6d1040017Ab0162bf00000100820008017Ab0162bf",
		INITVAL_1A => "0x000760006e0C4000D8000C8000E6000C27200067000420E6610E46b000690406109C000C2200D46f",
		INITVAL_1B => "0x0000000000000ff000ff00000000000000000000000000000000000000650006c000720006c00075",
		INITVAL_1C => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000",
		INITVAL_1D => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DIA0 => dmem_write_out(16), DIA1 => dmem_write_out(17),
		DIA2 => dmem_write_out(18), DIA3 => dmem_write_out(19),
		DIA4 => dmem_write_out(20), DIA5 => dmem_write_out(21),
		DIA6 => dmem_write_out(22), DIA7 => dmem_write_out(23),
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(16), DOA1 => dmem_data_read(17),
		DOA2 => dmem_data_read(18), DOA3 => dmem_data_read(19),
		DOA4 => dmem_data_read(20), DOA5 => dmem_data_read(21),
		DOA6 => dmem_data_read(22), DOA7 => dmem_data_read(23),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => dmem_addr(2), ADA4 => dmem_addr(3),
		ADA5 => dmem_addr(4), ADA6 => dmem_addr(5),
		ADA7 => dmem_addr(6), ADA8 => dmem_addr(7),
		ADA9 => dmem_addr(8), ADA10 => dmem_addr(9),
		ADA11 => dmem_addr(10), ADA12 => dmem_addr(11),
		ADA13 => dmem_addr(12),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_byte_we(2),
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(16), DOB1 => imem_data_out(17),
		DOB2 => imem_data_out(18), DOB3 => imem_data_out(19),
		DOB4 => imem_data_out(20), DOB5 => imem_data_out(21),
		DOB6 => imem_data_out(22), DOB7 => imem_data_out(23),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => imem_addr(2), ADB4 => imem_addr(3),
		ADB5 => imem_addr(4), ADB6 => imem_addr(5),
		ADB7 => imem_addr(6), ADB8 => imem_addr(7),
		ADB9 => imem_addr(8), ADB10 => imem_addr(9),
		ADB11 => imem_addr(10), ADB12 => imem_addr(11),
		ADB13 => imem_addr(12),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_3: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B=> "NORMAL", WRITEMODE_A => "NORMAL",
		GSR=> "DISABLED", RESETMODE=> "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A=> "NOREG",
		DATA_WIDTH_B=> 9, DATA_WIDTH_A=> 9,
		INITVAL_00 => "0x0489000018000000000015814048001180000025000240001406000028280001011E3c0183c06E3c",
		INITVAL_01 => "0x00018000000002500014048ac0000000000048000000000024000140600002828000030481414024",
		INITVAL_02 => "0x0202400624028300488c000140600000003048141002400010100000203000003048141402400000",
		INITVAL_03 => "0x06800000110581000015000000480006000002100480800000000000000300014000000001006000",
		INITVAL_04 => "0x0000000000000000000000000000000000011E270183407834078af0282711E00006ac0001000214",
		INITVAL_05 => "0x00000048260008f0040c0480004E0800400008af15Eaf15E2704E0315E000683c11E040000000000",
		INITVAL_06 => "0x14024048080002404808000a0048270068f11E8f11E140042614426144821048f0108f0280214414",
		INITVAL_07 => "0x12424048240000015Eaf15Eaf15Eaf15Eaf15Eaf04E2700003048141402400010050240480004810",
		INITVAL_08 => "0x01000020af01824118270068f11E8f11E8f004020108f0202c0200004C9204C1404C9211E1004C10",
		INITVAL_09 => "0x11E14000100000015E8f11E8f11E3002800000020001006010000000683c00010000af15Eaf04E02",
		INITVAL_0A => "0x00024048000683c15E1415Eaf04E8f00000000270068f11E2404E0311E8f11E140000011E00018af",
		INITVAL_0B => "0x15E00028000008f0683c11Eaf048af0480002824000140000011E8f15E00028000008f11Eaf15E24",
		INITVAL_0C => "0x000140500011E8f15E2415E8e0482404824048240482604E3104E0011Eaf048140000011E340788f",
		INITVAL_0D => "0x060100608f0000004800020280282800011000000008f1188f000100002500200028280008f11Eaf",
		INITVAL_0E => "0x04E0311E8f11E1604Caf028af000240001404800028280008f11Eaf000140500011E8f15Eaf00000",
		INITVAL_0F => "0x0042700400000af15E000608f0001015Eaf15Eaf15Eaf15E270000000208052010102e0521600012",
		INITVAL_10 => "0x15E8e04E0311E8f11E8f11E8f11E2602C26028020048e048000042700400000300008f0480c04802",
		INITVAL_11 => "0x0040004E0c15Eaf15Eaf15E02000af118af000270002715E08000300008f000080000c0048f0040c",
		INITVAL_12 => "0x11E8f11E8f11E8f11E0002024018240188f15E0c15E380002c0488f024240242402424024240040c",
		INITVAL_13 => "0x004020188e0040c0040000424000020040c00032118020642411E2702C24018260480204C2704E03",
		INITVAL_14 => "0x15E240001006000018340788f0480c0002407800018000000004E8e11C00000270040c0040004800",
		INITVAL_15 => "0x04C0c0008f0480002824018240188f11E140480c0480c11E24010af04E0811E8f11E8f11E8f11E24",
		INITVAL_16 => "0x0180011E140040c0002411E00018240000c00024010240188f0001611E140480c11E0c048140480c",
		INITVAL_17 => "0x11E300182411Eaf01800060000000c048080600c0002411E30018000008f004080008f0480c04824",
		INITVAL_18 => "0x15E100502411E100000011E8f11E0202C24018260480204Caf15E2715E270000000000010000608f",
		INITVAL_19 => "0x000720DA690A4000CC730CA6b00061040740E80015E0804E8f11E8f0000815Eaf010af04E8f11E8f",
		INITVAL_1A => "0x00065000690E4000D2000C2000E0000C66c00072000720D6760006f000630D6740C2000CC730CA6c",
		INITVAL_1B => "0x0000000000000ff000ff00000000000000000000000000000000000000650006c000650006500074",
		INITVAL_1C => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000",
		INITVAL_1D => "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000"
	)
	port map (
		DIA0 => dmem_write_out(24), DIA1 => dmem_write_out(25),
		DIA2 => dmem_write_out(26), DIA3 => dmem_write_out(27),
		DIA4 => dmem_write_out(28), DIA5 => dmem_write_out(29),
		DIA6 => dmem_write_out(30), DIA7 => dmem_write_out(31),
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(24), DOA1 => dmem_data_read(25),
		DOA2 => dmem_data_read(26), DOA3 => dmem_data_read(27),
		DOA4 => dmem_data_read(28), DOA5 => dmem_data_read(29),
		DOA6 => dmem_data_read(30), DOA7 => dmem_data_read(31),
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0', ADA2 => '0', 
		ADA3 => dmem_addr(2), ADA4 => dmem_addr(3),
		ADA5 => dmem_addr(4), ADA6 => dmem_addr(5),
		ADA7 => dmem_addr(6), ADA8 => dmem_addr(7),
		ADA9 => dmem_addr(8), ADA10 => dmem_addr(9),
		ADA11 => dmem_addr(10), ADA12 => dmem_addr(11),
		ADA13 => dmem_addr(12),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_byte_we(3),
		CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(24), DOB1 => imem_data_out(25),
		DOB2 => imem_data_out(26), DOB3 => imem_data_out(27),
		DOB4 => imem_data_out(28), DOB5 => imem_data_out(29),
		DOB6 => imem_data_out(30), DOB7 => imem_data_out(31),
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0', ADB2 => '0', 
		ADB3 => imem_addr(2), ADB4 => imem_addr(3),
		ADB5 => imem_addr(4), ADB6 => imem_addr(5),
		ADB7 => imem_addr(6), ADB8 => imem_addr(7),
		ADB9 => imem_addr(8), ADB10 => imem_addr(9),
		ADB11 => imem_addr(10), ADB12 => imem_addr(11),
		ADB13 => imem_addr(12),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

end Behavioral;
