library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package bootloader is
  type boot_block_type is array(0 to 511) of std_logic_vector(7 downto 0);

constant boot_block : boot_block_type := (
	x"00", x"00", x"00", x"00", x"21", x"40", x"00", x"00", 
	x"21", x"30", x"00", x"00", x"66", x"33", x"0a", x"3c", 
	x"3e", x"20", x"0b", x"3c", x"00", x"08", x"0c", x"3c", 
	x"01", x"00", x"0d", x"24", x"03", x"00", x"0e", x"24", 
	x"53", x"00", x"0f", x"24", x"0d", x"00", x"18", x"24", 
	x"21", x"c8", x"00", x"00", x"0d", x"0a", x"43", x"25", 
	x"21", x"ff", x"05", x"80", x"04", x"00", x"a7", x"30", 
	x"fd", x"ff", x"e0", x"14", x"00", x"00", x"00", x"00", 
	x"20", x"ff", x"03", x"a0", x"03", x"1a", x"03", x"00", 
	x"25", x"48", x"79", x"00", x"04", x"00", x"20", x"15", 
	x"00", x"00", x"00", x"00", x"ff", x"ff", x"19", x"24", 
	x"0c", x"00", x"00", x"08", x"32", x"63", x"63", x"25", 
	x"f3", x"ff", x"60", x"14", x"ff", x"00", x"05", x"24", 
	x"ff", x"ff", x"03", x"24", x"02", x"00", x"07", x"24", 
	x"1b", x"00", x"61", x"04", x"00", x"00", x"00", x"00", 
	x"00", x"48", x"02", x"40", x"24", x"c8", x"4c", x"00", 
	x"02", x"00", x"20", x"13", x"21", x"20", x"00", x"00", 
	x"ff", x"00", x"04", x"24", x"c3", x"cc", x"02", x"00", 
	x"ff", x"00", x"49", x"30", x"ff", x"00", x"39", x"33", 
	x"2a", x"48", x"29", x"03", x"03", x"00", x"20", x"11", 
	x"00", x"00", x"00", x"00", x"2c", x"00", x"00", x"08", 
	x"0f", x"00", x"84", x"38", x"f0", x"00", x"84", x"38", 
	x"11", x"ff", x"04", x"a0", x"21", x"ff", x"04", x"80", 
	x"01", x"00", x"99", x"30", x"ec", x"ff", x"20", x"13", 
	x"00", x"00", x"00", x"00", x"20", x"ff", x"04", x"80", 
	x"11", x"00", x"61", x"04", x"f6", x"ff", x"89", x"24", 
	x"05", x"00", x"8f", x"14", x"00", x"00", x"00", x"00", 
	x"21", x"10", x"00", x"00", x"21", x"18", x"00", x"00", 
	x"2c", x"00", x"00", x"08", x"03", x"22", x"06", x"00", 
	x"cf", x"ff", x"98", x"10", x"20", x"00", x"99", x"28", 
	x"df", x"ff", x"20", x"17", x"21", x"10", x"00", x"00", 
	x"21", x"ff", x"02", x"80", x"04", x"00", x"42", x"30", 
	x"fd", x"ff", x"40", x"14", x"00", x"00", x"00", x"00", 
	x"1c", x"00", x"00", x"08", x"20", x"ff", x"04", x"a0", 
	x"04", x"00", x"39", x"2d", x"05", x"00", x"20", x"13", 
	x"00", x"49", x"02", x"00", x"ff", x"00", x"05", x"24", 
	x"ff", x"ff", x"03", x"24", x"1e", x"00", x"00", x"08", 
	x"02", x"00", x"07", x"24", x"61", x"00", x"82", x"28", 
	x"03", x"00", x"40", x"14", x"d0", x"ff", x"82", x"24", 
	x"53", x"00", x"00", x"08", x"e0", x"ff", x"84", x"24", 
	x"41", x"00", x"99", x"28", x"03", x"00", x"20", x"17", 
	x"25", x"10", x"49", x"00", x"c9", x"ff", x"84", x"24", 
	x"25", x"10", x"89", x"00", x"01", x"00", x"63", x"24", 
	x"11", x"00", x"6d", x"14", x"f9", x"ff", x"59", x"24", 
	x"03", x"00", x"24", x"2f", x"09", x"00", x"80", x"10", 
	x"04", x"00", x"49", x"28", x"00", x"80", x"04", x"3c", 
	x"10", x"00", x"05", x"3c", x"24", x"e8", x"04", x"01", 
	x"21", x"f8", x"00", x"00", x"08", x"00", x"00", x"01", 
	x"25", x"e8", x"a5", x"03", x"1c", x"00", x"00", x"08", 
	x"21", x"10", x"00", x"00", x"fd", x"ff", x"20", x"11", 
	x"00", x"00", x"00", x"00", x"21", x"28", x"42", x"00", 
	x"61", x"00", x"00", x"08", x"05", x"00", x"a5", x"24", 
	x"04", x"00", x"6e", x"14", x"06", x"00", x"a9", x"28", 
	x"21", x"10", x"42", x"00", x"61", x"00", x"00", x"08", 
	x"21", x"38", x"e2", x"00", x"ae", x"ff", x"20", x"15", 
	x"00", x"00", x"00", x"00", x"06", x"00", x"65", x"14", 
	x"2a", x"c8", x"a3", x"00", x"02", x"00", x"00", x"15", 
	x"21", x"30", x"40", x"00", x"21", x"40", x"40", x"00", 
	x"1c", x"00", x"00", x"08", x"21", x"28", x"60", x"00", 
	x"a5", x"ff", x"20", x"13", x"01", x"00", x"64", x"30", 
	x"a3", x"ff", x"80", x"10", x"2a", x"48", x"67", x"00", 
	x"a1", x"ff", x"20", x"11", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"c2", x"a0", x"1c", x"00", x"00", x"08", 
	x"01", x"00", x"c6", x"24", x"00", x"00", x"00", x"00", 
	others => (others => '0')
    );

end bootloader;
