library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.font_block_pack.all;

package font8x16_xark is

constant font8x16_block : font16_block_type := (
		-- lines 1/1
		-- char 0x00='\0' 
		 0 =>	"00000000",	-- ........
		 1 =>	"00000000",	-- ........
		 2 =>	"00000000",	-- ........
		 3 =>	"00000000",	-- ........
		 4 =>	"00000000",	-- ........
		 5 =>	"00000000",	-- ........
		 6 =>	"00000000",	-- ........
		 7 =>	"00000000",	-- ........
		 8 =>	"00000000",	-- ........
		 9 =>	"00000000",	-- ........
		10 =>	"00000000",	-- ........
		11 =>	"00000000",	-- ........
		12 =>	"00000000",	-- ........
		13 =>	"00000000",	-- ........
		14 =>	"00000000",	-- ........
		15 =>	"00000000",	-- ........

		-- char 0x01='\x01
		16 =>	"00000000",	-- ........
		17 =>	"00000000",	-- ........
		18 =>	"00000000",	-- ........
		19 =>	"01111110",	-- .######.
		20 =>	"10000001",	-- #......#
		21 =>	"10100101",	-- #.#..#.#
		22 =>	"10000001",	-- #......#
		23 =>	"10000001",	-- #......#
		24 =>	"10111101",	-- #.####.#
		25 =>	"10011001",	-- #..##..#
		26 =>	"10000001",	-- #......#
		27 =>	"01111110",	-- .######.
		28 =>	"00000000",	-- ........
		29 =>	"00000000",	-- ........
		30 =>	"00000000",	-- ........
		31 =>	"00000000",	-- ........

		-- char 0x02='\x02
		32 =>	"00000000",	-- ........
		33 =>	"00000000",	-- ........
		34 =>	"00000000",	-- ........
		35 =>	"01111110",	-- .######.
		36 =>	"11111111",	-- ########
		37 =>	"11011011",	-- ##.##.##
		38 =>	"11111111",	-- ########
		39 =>	"11111111",	-- ########
		40 =>	"11000011",	-- ##....##
		41 =>	"11100111",	-- ###..###
		42 =>	"11111111",	-- ########
		43 =>	"01111110",	-- .######.
		44 =>	"00000000",	-- ........
		45 =>	"00000000",	-- ........
		46 =>	"00000000",	-- ........
		47 =>	"00000000",	-- ........

		-- char 0x03='\x03
		48 =>	"00000000",	-- ........
		49 =>	"00000000",	-- ........
		50 =>	"00000000",	-- ........
		51 =>	"00000000",	-- ........
		52 =>	"01101100",	-- .##.##..
		53 =>	"11111110",	-- #######.
		54 =>	"11111110",	-- #######.
		55 =>	"11111110",	-- #######.
		56 =>	"11111110",	-- #######.
		57 =>	"01111100",	-- .#####..
		58 =>	"00111000",	-- ..###...
		59 =>	"00010000",	-- ...#....
		60 =>	"00000000",	-- ........
		61 =>	"00000000",	-- ........
		62 =>	"00000000",	-- ........
		63 =>	"00000000",	-- ........

		-- char 0x04='\x04
		64 =>	"00000000",	-- ........
		65 =>	"00000000",	-- ........
		66 =>	"00000000",	-- ........
		67 =>	"00000000",	-- ........
		68 =>	"00010000",	-- ...#....
		69 =>	"00111000",	-- ..###...
		70 =>	"01111100",	-- .#####..
		71 =>	"11111110",	-- #######.
		72 =>	"01111100",	-- .#####..
		73 =>	"00111000",	-- ..###...
		74 =>	"00010000",	-- ...#....
		75 =>	"00000000",	-- ........
		76 =>	"00000000",	-- ........
		77 =>	"00000000",	-- ........
		78 =>	"00000000",	-- ........
		79 =>	"00000000",	-- ........

		-- char 0x05='\x05
		80 =>	"00000000",	-- ........
		81 =>	"00000000",	-- ........
		82 =>	"00000000",	-- ........
		83 =>	"00011000",	-- ...##...
		84 =>	"00111100",	-- ..####..
		85 =>	"00111100",	-- ..####..
		86 =>	"11100111",	-- ###..###
		87 =>	"11100111",	-- ###..###
		88 =>	"11100111",	-- ###..###
		89 =>	"00011000",	-- ...##...
		90 =>	"00011000",	-- ...##...
		91 =>	"00111100",	-- ..####..
		92 =>	"00000000",	-- ........
		93 =>	"00000000",	-- ........
		94 =>	"00000000",	-- ........
		95 =>	"00000000",	-- ........

		-- char 0x06='\x06
		96 =>	"00000000",	-- ........
		97 =>	"00000000",	-- ........
		98 =>	"00000000",	-- ........
		99 =>	"00011000",	-- ...##...
		100 =>	"00111100",	-- ..####..
		101 =>	"01111110",	-- .######.
		102 =>	"11111111",	-- ########
		103 =>	"11111111",	-- ########
		104 =>	"01111110",	-- .######.
		105 =>	"00011000",	-- ...##...
		106 =>	"00011000",	-- ...##...
		107 =>	"00111100",	-- ..####..
		108 =>	"00000000",	-- ........
		109 =>	"00000000",	-- ........
		110 =>	"00000000",	-- ........
		111 =>	"00000000",	-- ........

		-- char 0x07='\a' 
		112 =>	"00000000",	-- ........
		113 =>	"00000000",	-- ........
		114 =>	"00000000",	-- ........
		115 =>	"00000000",	-- ........
		116 =>	"00000000",	-- ........
		117 =>	"00000000",	-- ........
		118 =>	"00011000",	-- ...##...
		119 =>	"00111100",	-- ..####..
		120 =>	"00111100",	-- ..####..
		121 =>	"00011000",	-- ...##...
		122 =>	"00000000",	-- ........
		123 =>	"00000000",	-- ........
		124 =>	"00000000",	-- ........
		125 =>	"00000000",	-- ........
		126 =>	"00000000",	-- ........
		127 =>	"00000000",	-- ........

		-- char 0x08='\b' 
		128 =>	"11111111",	-- ########
		129 =>	"11111111",	-- ########
		130 =>	"11111111",	-- ########
		131 =>	"11111111",	-- ########
		132 =>	"11111111",	-- ########
		133 =>	"11111111",	-- ########
		134 =>	"11100111",	-- ###..###
		135 =>	"11000011",	-- ##....##
		136 =>	"11000011",	-- ##....##
		137 =>	"11100111",	-- ###..###
		138 =>	"11111111",	-- ########
		139 =>	"11111111",	-- ########
		140 =>	"11111111",	-- ########
		141 =>	"11111111",	-- ########
		142 =>	"11111111",	-- ########
		143 =>	"11111111",	-- ########

		-- char 0x09='\t' 
		144 =>	"00000000",	-- ........
		145 =>	"00000000",	-- ........
		146 =>	"00000000",	-- ........
		147 =>	"00000000",	-- ........
		148 =>	"00000000",	-- ........
		149 =>	"00111100",	-- ..####..
		150 =>	"01100110",	-- .##..##.
		151 =>	"01000010",	-- .#....#.
		152 =>	"01000010",	-- .#....#.
		153 =>	"01100110",	-- .##..##.
		154 =>	"00111100",	-- ..####..
		155 =>	"00000000",	-- ........
		156 =>	"00000000",	-- ........
		157 =>	"00000000",	-- ........
		158 =>	"00000000",	-- ........
		159 =>	"00000000",	-- ........

		-- char 0x0a='\n' 
		160 =>	"00000000",	-- ........
		161 =>	"11111111",	-- ########
		162 =>	"11111111",	-- ########
		163 =>	"11111111",	-- ########
		164 =>	"11111111",	-- ########
		165 =>	"11000011",	-- ##....##
		166 =>	"10011001",	-- #..##..#
		167 =>	"10111101",	-- #.####.#
		168 =>	"10111101",	-- #.####.#
		169 =>	"10011001",	-- #..##..#
		170 =>	"11000011",	-- ##....##
		171 =>	"11111111",	-- ########
		172 =>	"11111111",	-- ########
		173 =>	"11111111",	-- ########
		174 =>	"11111111",	-- ########
		175 =>	"00000000",	-- ........

		-- char 0x0b='\v' 
		176 =>	"00000000",	-- ........
		177 =>	"00000000",	-- ........
		178 =>	"00000000",	-- ........
		179 =>	"00011110",	-- ...####.
		180 =>	"00001110",	-- ....###.
		181 =>	"00011010",	-- ...##.#.
		182 =>	"00110010",	-- ..##..#.
		183 =>	"01111000",	-- .####...
		184 =>	"11001100",	-- ##..##..
		185 =>	"11001100",	-- ##..##..
		186 =>	"11001100",	-- ##..##..
		187 =>	"01111000",	-- .####...
		188 =>	"00000000",	-- ........
		189 =>	"00000000",	-- ........
		190 =>	"00000000",	-- ........
		191 =>	"00000000",	-- ........

		-- char 0x0c='\f' 
		192 =>	"00000000",	-- ........
		193 =>	"00000000",	-- ........
		194 =>	"00000000",	-- ........
		195 =>	"00111100",	-- ..####..
		196 =>	"01100110",	-- .##..##.
		197 =>	"01100110",	-- .##..##.
		198 =>	"01100110",	-- .##..##.
		199 =>	"00111100",	-- ..####..
		200 =>	"00011000",	-- ...##...
		201 =>	"01111110",	-- .######.
		202 =>	"00011000",	-- ...##...
		203 =>	"00011000",	-- ...##...
		204 =>	"00000000",	-- ........
		205 =>	"00000000",	-- ........
		206 =>	"00000000",	-- ........
		207 =>	"00000000",	-- ........

		-- char 0x0d='\r' 
		208 =>	"00000000",	-- ........
		209 =>	"00000000",	-- ........
		210 =>	"00000000",	-- ........
		211 =>	"00111111",	-- ..######
		212 =>	"00110011",	-- ..##..##
		213 =>	"00111111",	-- ..######
		214 =>	"00110000",	-- ..##....
		215 =>	"00110000",	-- ..##....
		216 =>	"00110000",	-- ..##....
		217 =>	"01110000",	-- .###....
		218 =>	"11110000",	-- ####....
		219 =>	"11100000",	-- ###.....
		220 =>	"00000000",	-- ........
		221 =>	"00000000",	-- ........
		222 =>	"00000000",	-- ........
		223 =>	"00000000",	-- ........

		-- char 0x0e='\x0e
		224 =>	"00000000",	-- ........
		225 =>	"00000000",	-- ........
		226 =>	"00000000",	-- ........
		227 =>	"01111111",	-- .#######
		228 =>	"01100011",	-- .##...##
		229 =>	"01111111",	-- .#######
		230 =>	"01100011",	-- .##...##
		231 =>	"01100011",	-- .##...##
		232 =>	"01100011",	-- .##...##
		233 =>	"01100111",	-- .##..###
		234 =>	"11100111",	-- ###..###
		235 =>	"11100110",	-- ###..##.
		236 =>	"11000000",	-- ##......
		237 =>	"00000000",	-- ........
		238 =>	"00000000",	-- ........
		239 =>	"00000000",	-- ........

		-- char 0x0f='\x0f
		240 =>	"00000000",	-- ........
		241 =>	"00000000",	-- ........
		242 =>	"00000000",	-- ........
		243 =>	"00011000",	-- ...##...
		244 =>	"00011000",	-- ...##...
		245 =>	"11011011",	-- ##.##.##
		246 =>	"00111100",	-- ..####..
		247 =>	"11100111",	-- ###..###
		248 =>	"00111100",	-- ..####..
		249 =>	"11011011",	-- ##.##.##
		250 =>	"00011000",	-- ...##...
		251 =>	"00011000",	-- ...##...
		252 =>	"00000000",	-- ........
		253 =>	"00000000",	-- ........
		254 =>	"00000000",	-- ........
		255 =>	"00000000",	-- ........

		-- char 0x10='\x10
		256 =>	"00000000",	-- ........
		257 =>	"00000000",	-- ........
		258 =>	"00000000",	-- ........
		259 =>	"10000000",	-- #.......
		260 =>	"11000000",	-- ##......
		261 =>	"11100000",	-- ###.....
		262 =>	"11111000",	-- #####...
		263 =>	"11111110",	-- #######.
		264 =>	"11111000",	-- #####...
		265 =>	"11100000",	-- ###.....
		266 =>	"11000000",	-- ##......
		267 =>	"10000000",	-- #.......
		268 =>	"00000000",	-- ........
		269 =>	"00000000",	-- ........
		270 =>	"00000000",	-- ........
		271 =>	"00000000",	-- ........

		-- char 0x11='\x11
		272 =>	"00000000",	-- ........
		273 =>	"00000000",	-- ........
		274 =>	"00000000",	-- ........
		275 =>	"00000010",	-- ......#.
		276 =>	"00000110",	-- .....##.
		277 =>	"00001110",	-- ....###.
		278 =>	"00111110",	-- ..#####.
		279 =>	"11111110",	-- #######.
		280 =>	"00111110",	-- ..#####.
		281 =>	"00001110",	-- ....###.
		282 =>	"00000110",	-- .....##.
		283 =>	"00000010",	-- ......#.
		284 =>	"00000000",	-- ........
		285 =>	"00000000",	-- ........
		286 =>	"00000000",	-- ........
		287 =>	"00000000",	-- ........

		-- char 0x12='\x12
		288 =>	"00000000",	-- ........
		289 =>	"00000000",	-- ........
		290 =>	"00000000",	-- ........
		291 =>	"00011000",	-- ...##...
		292 =>	"00111100",	-- ..####..
		293 =>	"01111110",	-- .######.
		294 =>	"00011000",	-- ...##...
		295 =>	"00011000",	-- ...##...
		296 =>	"00011000",	-- ...##...
		297 =>	"01111110",	-- .######.
		298 =>	"00111100",	-- ..####..
		299 =>	"00011000",	-- ...##...
		300 =>	"00000000",	-- ........
		301 =>	"00000000",	-- ........
		302 =>	"00000000",	-- ........
		303 =>	"00000000",	-- ........

		-- char 0x13='\x13
		304 =>	"00000000",	-- ........
		305 =>	"00000000",	-- ........
		306 =>	"00000000",	-- ........
		307 =>	"01100110",	-- .##..##.
		308 =>	"01100110",	-- .##..##.
		309 =>	"01100110",	-- .##..##.
		310 =>	"01100110",	-- .##..##.
		311 =>	"01100110",	-- .##..##.
		312 =>	"01100110",	-- .##..##.
		313 =>	"00000000",	-- ........
		314 =>	"01100110",	-- .##..##.
		315 =>	"01100110",	-- .##..##.
		316 =>	"00000000",	-- ........
		317 =>	"00000000",	-- ........
		318 =>	"00000000",	-- ........
		319 =>	"00000000",	-- ........

		-- char 0x14='\x14
		320 =>	"00000000",	-- ........
		321 =>	"00000000",	-- ........
		322 =>	"00000000",	-- ........
		323 =>	"01111111",	-- .#######
		324 =>	"11011011",	-- ##.##.##
		325 =>	"11011011",	-- ##.##.##
		326 =>	"11011011",	-- ##.##.##
		327 =>	"01111011",	-- .####.##
		328 =>	"00011011",	-- ...##.##
		329 =>	"00011011",	-- ...##.##
		330 =>	"00011011",	-- ...##.##
		331 =>	"00011011",	-- ...##.##
		332 =>	"00000000",	-- ........
		333 =>	"00000000",	-- ........
		334 =>	"00000000",	-- ........
		335 =>	"00000000",	-- ........

		-- char 0x15='\x15
		336 =>	"00000000",	-- ........
		337 =>	"00000000",	-- ........
		338 =>	"01111100",	-- .#####..
		339 =>	"11000110",	-- ##...##.
		340 =>	"01100000",	-- .##.....
		341 =>	"00111000",	-- ..###...
		342 =>	"01101100",	-- .##.##..
		343 =>	"11000110",	-- ##...##.
		344 =>	"11000110",	-- ##...##.
		345 =>	"01101100",	-- .##.##..
		346 =>	"00111000",	-- ..###...
		347 =>	"00001100",	-- ....##..
		348 =>	"11000110",	-- ##...##.
		349 =>	"01111100",	-- .#####..
		350 =>	"00000000",	-- ........
		351 =>	"00000000",	-- ........

		-- char 0x16='\x16
		352 =>	"00000000",	-- ........
		353 =>	"00000000",	-- ........
		354 =>	"00000000",	-- ........
		355 =>	"00000000",	-- ........
		356 =>	"00000000",	-- ........
		357 =>	"00000000",	-- ........
		358 =>	"00000000",	-- ........
		359 =>	"00000000",	-- ........
		360 =>	"00000000",	-- ........
		361 =>	"11111110",	-- #######.
		362 =>	"11111110",	-- #######.
		363 =>	"11111110",	-- #######.
		364 =>	"00000000",	-- ........
		365 =>	"00000000",	-- ........
		366 =>	"00000000",	-- ........
		367 =>	"00000000",	-- ........

		-- char 0x17='\x17
		368 =>	"00000000",	-- ........
		369 =>	"00000000",	-- ........
		370 =>	"00000000",	-- ........
		371 =>	"00011000",	-- ...##...
		372 =>	"00111100",	-- ..####..
		373 =>	"01111110",	-- .######.
		374 =>	"00011000",	-- ...##...
		375 =>	"00011000",	-- ...##...
		376 =>	"00011000",	-- ...##...
		377 =>	"01111110",	-- .######.
		378 =>	"00111100",	-- ..####..
		379 =>	"00011000",	-- ...##...
		380 =>	"01111110",	-- .######.
		381 =>	"00000000",	-- ........
		382 =>	"00000000",	-- ........
		383 =>	"00000000",	-- ........

		-- char 0x18='\x18
		384 =>	"00000000",	-- ........
		385 =>	"00000000",	-- ........
		386 =>	"00000000",	-- ........
		387 =>	"00011000",	-- ...##...
		388 =>	"00111100",	-- ..####..
		389 =>	"01111110",	-- .######.
		390 =>	"00011000",	-- ...##...
		391 =>	"00011000",	-- ...##...
		392 =>	"00011000",	-- ...##...
		393 =>	"00011000",	-- ...##...
		394 =>	"00011000",	-- ...##...
		395 =>	"00011000",	-- ...##...
		396 =>	"00000000",	-- ........
		397 =>	"00000000",	-- ........
		398 =>	"00000000",	-- ........
		399 =>	"00000000",	-- ........

		-- char 0x19='\x19
		400 =>	"00000000",	-- ........
		401 =>	"00000000",	-- ........
		402 =>	"00000000",	-- ........
		403 =>	"00011000",	-- ...##...
		404 =>	"00011000",	-- ...##...
		405 =>	"00011000",	-- ...##...
		406 =>	"00011000",	-- ...##...
		407 =>	"00011000",	-- ...##...
		408 =>	"00011000",	-- ...##...
		409 =>	"01111110",	-- .######.
		410 =>	"00111100",	-- ..####..
		411 =>	"00011000",	-- ...##...
		412 =>	"00000000",	-- ........
		413 =>	"00000000",	-- ........
		414 =>	"00000000",	-- ........
		415 =>	"00000000",	-- ........

		-- char 0x1a='\x1a
		416 =>	"00000000",	-- ........
		417 =>	"00000000",	-- ........
		418 =>	"00000000",	-- ........
		419 =>	"00000000",	-- ........
		420 =>	"00000000",	-- ........
		421 =>	"00011000",	-- ...##...
		422 =>	"00001100",	-- ....##..
		423 =>	"11111110",	-- #######.
		424 =>	"00001100",	-- ....##..
		425 =>	"00011000",	-- ...##...
		426 =>	"00000000",	-- ........
		427 =>	"00000000",	-- ........
		428 =>	"00000000",	-- ........
		429 =>	"00000000",	-- ........
		430 =>	"00000000",	-- ........
		431 =>	"00000000",	-- ........

		-- char 0x1b='\x1b
		432 =>	"00000000",	-- ........
		433 =>	"00000000",	-- ........
		434 =>	"00000000",	-- ........
		435 =>	"00000000",	-- ........
		436 =>	"00000000",	-- ........
		437 =>	"00110000",	-- ..##....
		438 =>	"01100000",	-- .##.....
		439 =>	"11111110",	-- #######.
		440 =>	"01100000",	-- .##.....
		441 =>	"00110000",	-- ..##....
		442 =>	"00000000",	-- ........
		443 =>	"00000000",	-- ........
		444 =>	"00000000",	-- ........
		445 =>	"00000000",	-- ........
		446 =>	"00000000",	-- ........
		447 =>	"00000000",	-- ........

		-- char 0x1c='\x1c
		448 =>	"00000000",	-- ........
		449 =>	"00000000",	-- ........
		450 =>	"00000000",	-- ........
		451 =>	"00000000",	-- ........
		452 =>	"00000000",	-- ........
		453 =>	"00000000",	-- ........
		454 =>	"11000000",	-- ##......
		455 =>	"11000000",	-- ##......
		456 =>	"11000000",	-- ##......
		457 =>	"11111110",	-- #######.
		458 =>	"00000000",	-- ........
		459 =>	"00000000",	-- ........
		460 =>	"00000000",	-- ........
		461 =>	"00000000",	-- ........
		462 =>	"00000000",	-- ........
		463 =>	"00000000",	-- ........

		-- char 0x1d='\x1d
		464 =>	"00000000",	-- ........
		465 =>	"00000000",	-- ........
		466 =>	"00000000",	-- ........
		467 =>	"00000000",	-- ........
		468 =>	"00000000",	-- ........
		469 =>	"00101000",	-- ..#.#...
		470 =>	"01101100",	-- .##.##..
		471 =>	"11111110",	-- #######.
		472 =>	"01101100",	-- .##.##..
		473 =>	"00101000",	-- ..#.#...
		474 =>	"00000000",	-- ........
		475 =>	"00000000",	-- ........
		476 =>	"00000000",	-- ........
		477 =>	"00000000",	-- ........
		478 =>	"00000000",	-- ........
		479 =>	"00000000",	-- ........

		-- char 0x1e='\x1e
		480 =>	"00000000",	-- ........
		481 =>	"00000000",	-- ........
		482 =>	"00000000",	-- ........
		483 =>	"00000000",	-- ........
		484 =>	"00010000",	-- ...#....
		485 =>	"00111000",	-- ..###...
		486 =>	"00111000",	-- ..###...
		487 =>	"01111100",	-- .#####..
		488 =>	"01111100",	-- .#####..
		489 =>	"11111110",	-- #######.
		490 =>	"11111110",	-- #######.
		491 =>	"00000000",	-- ........
		492 =>	"00000000",	-- ........
		493 =>	"00000000",	-- ........
		494 =>	"00000000",	-- ........
		495 =>	"00000000",	-- ........

		-- char 0x1f='\x1f
		496 =>	"00000000",	-- ........
		497 =>	"00000000",	-- ........
		498 =>	"00000000",	-- ........
		499 =>	"00000000",	-- ........
		500 =>	"11111110",	-- #######.
		501 =>	"11111110",	-- #######.
		502 =>	"01111100",	-- .#####..
		503 =>	"01111100",	-- .#####..
		504 =>	"00111000",	-- ..###...
		505 =>	"00111000",	-- ..###...
		506 =>	"00010000",	-- ...#....
		507 =>	"00000000",	-- ........
		508 =>	"00000000",	-- ........
		509 =>	"00000000",	-- ........
		510 =>	"00000000",	-- ........
		511 =>	"00000000",	-- ........

		-- char 0x20=' '  
		512 =>	"00000000",	-- ........
		513 =>	"00000000",	-- ........
		514 =>	"00000000",	-- ........
		515 =>	"00000000",	-- ........
		516 =>	"00000000",	-- ........
		517 =>	"00000000",	-- ........
		518 =>	"00000000",	-- ........
		519 =>	"00000000",	-- ........
		520 =>	"00000000",	-- ........
		521 =>	"00000000",	-- ........
		522 =>	"00000000",	-- ........
		523 =>	"00000000",	-- ........
		524 =>	"00000000",	-- ........
		525 =>	"00000000",	-- ........
		526 =>	"00000000",	-- ........
		527 =>	"00000000",	-- ........

		-- char 0x21='!'  
		528 =>	"00000000",	-- ........
		529 =>	"00000000",	-- ........
		530 =>	"00000000",	-- ........
		531 =>	"00011000",	-- ...##...
		532 =>	"00111100",	-- ..####..
		533 =>	"00111100",	-- ..####..
		534 =>	"00111100",	-- ..####..
		535 =>	"00011000",	-- ...##...
		536 =>	"00011000",	-- ...##...
		537 =>	"00000000",	-- ........
		538 =>	"00011000",	-- ...##...
		539 =>	"00011000",	-- ...##...
		540 =>	"00000000",	-- ........
		541 =>	"00000000",	-- ........
		542 =>	"00000000",	-- ........
		543 =>	"00000000",	-- ........

		-- char 0x22='\'' 
		544 =>	"00000000",	-- ........
		545 =>	"00000000",	-- ........
		546 =>	"01100110",	-- .##..##.
		547 =>	"01100110",	-- .##..##.
		548 =>	"01100110",	-- .##..##.
		549 =>	"00100100",	-- ..#..#..
		550 =>	"00000000",	-- ........
		551 =>	"00000000",	-- ........
		552 =>	"00000000",	-- ........
		553 =>	"00000000",	-- ........
		554 =>	"00000000",	-- ........
		555 =>	"00000000",	-- ........
		556 =>	"00000000",	-- ........
		557 =>	"00000000",	-- ........
		558 =>	"00000000",	-- ........
		559 =>	"00000000",	-- ........

		-- char 0x23='#'  
		560 =>	"00000000",	-- ........
		561 =>	"00000000",	-- ........
		562 =>	"00000000",	-- ........
		563 =>	"01101100",	-- .##.##..
		564 =>	"01101100",	-- .##.##..
		565 =>	"11111110",	-- #######.
		566 =>	"01101100",	-- .##.##..
		567 =>	"01101100",	-- .##.##..
		568 =>	"01101100",	-- .##.##..
		569 =>	"11111110",	-- #######.
		570 =>	"01101100",	-- .##.##..
		571 =>	"01101100",	-- .##.##..
		572 =>	"00000000",	-- ........
		573 =>	"00000000",	-- ........
		574 =>	"00000000",	-- ........
		575 =>	"00000000",	-- ........

		-- char 0x24='$'  
		576 =>	"00000000",	-- ........
		577 =>	"00011000",	-- ...##...
		578 =>	"00011000",	-- ...##...
		579 =>	"01111100",	-- .#####..
		580 =>	"11000110",	-- ##...##.
		581 =>	"11000010",	-- ##....#.
		582 =>	"11000000",	-- ##......
		583 =>	"01111100",	-- .#####..
		584 =>	"00000110",	-- .....##.
		585 =>	"10000110",	-- #....##.
		586 =>	"11000110",	-- ##...##.
		587 =>	"01111100",	-- .#####..
		588 =>	"00011000",	-- ...##...
		589 =>	"00011000",	-- ...##...
		590 =>	"00000000",	-- ........
		591 =>	"00000000",	-- ........

		-- char 0x25='%'  
		592 =>	"00000000",	-- ........
		593 =>	"00000000",	-- ........
		594 =>	"00000000",	-- ........
		595 =>	"00000000",	-- ........
		596 =>	"00000000",	-- ........
		597 =>	"11000010",	-- ##....#.
		598 =>	"11000110",	-- ##...##.
		599 =>	"00001100",	-- ....##..
		600 =>	"00011000",	-- ...##...
		601 =>	"00110000",	-- ..##....
		602 =>	"01100110",	-- .##..##.
		603 =>	"11000110",	-- ##...##.
		604 =>	"00000000",	-- ........
		605 =>	"00000000",	-- ........
		606 =>	"00000000",	-- ........
		607 =>	"00000000",	-- ........

		-- char 0x26='&'  
		608 =>	"00000000",	-- ........
		609 =>	"00000000",	-- ........
		610 =>	"00000000",	-- ........
		611 =>	"00111000",	-- ..###...
		612 =>	"01101100",	-- .##.##..
		613 =>	"01101100",	-- .##.##..
		614 =>	"00111000",	-- ..###...
		615 =>	"01110110",	-- .###.##.
		616 =>	"11011100",	-- ##.###..
		617 =>	"11001100",	-- ##..##..
		618 =>	"11001100",	-- ##..##..
		619 =>	"01110110",	-- .###.##.
		620 =>	"00000000",	-- ........
		621 =>	"00000000",	-- ........
		622 =>	"00000000",	-- ........
		623 =>	"00000000",	-- ........

		-- char 0x27='\"' 
		624 =>	"00000000",	-- ........
		625 =>	"00000000",	-- ........
		626 =>	"00110000",	-- ..##....
		627 =>	"00110000",	-- ..##....
		628 =>	"00110000",	-- ..##....
		629 =>	"01100000",	-- .##.....
		630 =>	"00000000",	-- ........
		631 =>	"00000000",	-- ........
		632 =>	"00000000",	-- ........
		633 =>	"00000000",	-- ........
		634 =>	"00000000",	-- ........
		635 =>	"00000000",	-- ........
		636 =>	"00000000",	-- ........
		637 =>	"00000000",	-- ........
		638 =>	"00000000",	-- ........
		639 =>	"00000000",	-- ........

		-- char 0x28='('  
		640 =>	"00000000",	-- ........
		641 =>	"00000000",	-- ........
		642 =>	"00000000",	-- ........
		643 =>	"00001100",	-- ....##..
		644 =>	"00011000",	-- ...##...
		645 =>	"00110000",	-- ..##....
		646 =>	"00110000",	-- ..##....
		647 =>	"00110000",	-- ..##....
		648 =>	"00110000",	-- ..##....
		649 =>	"00110000",	-- ..##....
		650 =>	"00011000",	-- ...##...
		651 =>	"00001100",	-- ....##..
		652 =>	"00000000",	-- ........
		653 =>	"00000000",	-- ........
		654 =>	"00000000",	-- ........
		655 =>	"00000000",	-- ........

		-- char 0x29=')'  
		656 =>	"00000000",	-- ........
		657 =>	"00000000",	-- ........
		658 =>	"00000000",	-- ........
		659 =>	"00110000",	-- ..##....
		660 =>	"00011000",	-- ...##...
		661 =>	"00001100",	-- ....##..
		662 =>	"00001100",	-- ....##..
		663 =>	"00001100",	-- ....##..
		664 =>	"00001100",	-- ....##..
		665 =>	"00001100",	-- ....##..
		666 =>	"00011000",	-- ...##...
		667 =>	"00110000",	-- ..##....
		668 =>	"00000000",	-- ........
		669 =>	"00000000",	-- ........
		670 =>	"00000000",	-- ........
		671 =>	"00000000",	-- ........

		-- char 0x2a='*'  
		672 =>	"00000000",	-- ........
		673 =>	"00000000",	-- ........
		674 =>	"00000000",	-- ........
		675 =>	"00000000",	-- ........
		676 =>	"00000000",	-- ........
		677 =>	"01100110",	-- .##..##.
		678 =>	"00111100",	-- ..####..
		679 =>	"11111111",	-- ########
		680 =>	"00111100",	-- ..####..
		681 =>	"01100110",	-- .##..##.
		682 =>	"00000000",	-- ........
		683 =>	"00000000",	-- ........
		684 =>	"00000000",	-- ........
		685 =>	"00000000",	-- ........
		686 =>	"00000000",	-- ........
		687 =>	"00000000",	-- ........

		-- char 0x2b='+'  
		688 =>	"00000000",	-- ........
		689 =>	"00000000",	-- ........
		690 =>	"00000000",	-- ........
		691 =>	"00000000",	-- ........
		692 =>	"00000000",	-- ........
		693 =>	"00011000",	-- ...##...
		694 =>	"00011000",	-- ...##...
		695 =>	"01111110",	-- .######.
		696 =>	"00011000",	-- ...##...
		697 =>	"00011000",	-- ...##...
		698 =>	"00000000",	-- ........
		699 =>	"00000000",	-- ........
		700 =>	"00000000",	-- ........
		701 =>	"00000000",	-- ........
		702 =>	"00000000",	-- ........
		703 =>	"00000000",	-- ........

		-- char 0x2c=','  
		704 =>	"00000000",	-- ........
		705 =>	"00000000",	-- ........
		706 =>	"00000000",	-- ........
		707 =>	"00000000",	-- ........
		708 =>	"00000000",	-- ........
		709 =>	"00000000",	-- ........
		710 =>	"00000000",	-- ........
		711 =>	"00000000",	-- ........
		712 =>	"00000000",	-- ........
		713 =>	"00011000",	-- ...##...
		714 =>	"00011000",	-- ...##...
		715 =>	"00011000",	-- ...##...
		716 =>	"00110000",	-- ..##....
		717 =>	"00000000",	-- ........
		718 =>	"00000000",	-- ........
		719 =>	"00000000",	-- ........

		-- char 0x2d='-'  
		720 =>	"00000000",	-- ........
		721 =>	"00000000",	-- ........
		722 =>	"00000000",	-- ........
		723 =>	"00000000",	-- ........
		724 =>	"00000000",	-- ........
		725 =>	"00000000",	-- ........
		726 =>	"00000000",	-- ........
		727 =>	"11111110",	-- #######.
		728 =>	"00000000",	-- ........
		729 =>	"00000000",	-- ........
		730 =>	"00000000",	-- ........
		731 =>	"00000000",	-- ........
		732 =>	"00000000",	-- ........
		733 =>	"00000000",	-- ........
		734 =>	"00000000",	-- ........
		735 =>	"00000000",	-- ........

		-- char 0x2e='.'  
		736 =>	"00000000",	-- ........
		737 =>	"00000000",	-- ........
		738 =>	"00000000",	-- ........
		739 =>	"00000000",	-- ........
		740 =>	"00000000",	-- ........
		741 =>	"00000000",	-- ........
		742 =>	"00000000",	-- ........
		743 =>	"00000000",	-- ........
		744 =>	"00000000",	-- ........
		745 =>	"00000000",	-- ........
		746 =>	"00011000",	-- ...##...
		747 =>	"00011000",	-- ...##...
		748 =>	"00000000",	-- ........
		749 =>	"00000000",	-- ........
		750 =>	"00000000",	-- ........
		751 =>	"00000000",	-- ........

		-- char 0x2f='/'  
		752 =>	"00000000",	-- ........
		753 =>	"00000000",	-- ........
		754 =>	"00000000",	-- ........
		755 =>	"00000010",	-- ......#.
		756 =>	"00000110",	-- .....##.
		757 =>	"00001100",	-- ....##..
		758 =>	"00011000",	-- ...##...
		759 =>	"00110000",	-- ..##....
		760 =>	"01100000",	-- .##.....
		761 =>	"11000000",	-- ##......
		762 =>	"10000000",	-- #.......
		763 =>	"00000000",	-- ........
		764 =>	"00000000",	-- ........
		765 =>	"00000000",	-- ........
		766 =>	"00000000",	-- ........
		767 =>	"00000000",	-- ........

		-- char 0x30='0'  
		768 =>	"00000000",	-- ........
		769 =>	"00000000",	-- ........
		770 =>	"00000000",	-- ........
		771 =>	"01111100",	-- .#####..
		772 =>	"11000110",	-- ##...##.
		773 =>	"11001110",	-- ##..###.
		774 =>	"11011110",	-- ##.####.
		775 =>	"11110110",	-- ####.##.
		776 =>	"11100110",	-- ###..##.
		777 =>	"11000110",	-- ##...##.
		778 =>	"11000110",	-- ##...##.
		779 =>	"01111100",	-- .#####..
		780 =>	"00000000",	-- ........
		781 =>	"00000000",	-- ........
		782 =>	"00000000",	-- ........
		783 =>	"00000000",	-- ........

		-- char 0x31='1'  
		784 =>	"00000000",	-- ........
		785 =>	"00000000",	-- ........
		786 =>	"00000000",	-- ........
		787 =>	"00011000",	-- ...##...
		788 =>	"00111000",	-- ..###...
		789 =>	"01111000",	-- .####...
		790 =>	"00011000",	-- ...##...
		791 =>	"00011000",	-- ...##...
		792 =>	"00011000",	-- ...##...
		793 =>	"00011000",	-- ...##...
		794 =>	"00011000",	-- ...##...
		795 =>	"01111110",	-- .######.
		796 =>	"00000000",	-- ........
		797 =>	"00000000",	-- ........
		798 =>	"00000000",	-- ........
		799 =>	"00000000",	-- ........

		-- char 0x32='2'  
		800 =>	"00000000",	-- ........
		801 =>	"00000000",	-- ........
		802 =>	"00000000",	-- ........
		803 =>	"01111100",	-- .#####..
		804 =>	"11000110",	-- ##...##.
		805 =>	"00000110",	-- .....##.
		806 =>	"00001100",	-- ....##..
		807 =>	"00011000",	-- ...##...
		808 =>	"00110000",	-- ..##....
		809 =>	"01100000",	-- .##.....
		810 =>	"11000110",	-- ##...##.
		811 =>	"11111110",	-- #######.
		812 =>	"00000000",	-- ........
		813 =>	"00000000",	-- ........
		814 =>	"00000000",	-- ........
		815 =>	"00000000",	-- ........

		-- char 0x33='3'  
		816 =>	"00000000",	-- ........
		817 =>	"00000000",	-- ........
		818 =>	"00000000",	-- ........
		819 =>	"01111100",	-- .#####..
		820 =>	"11000110",	-- ##...##.
		821 =>	"00000110",	-- .....##.
		822 =>	"00000110",	-- .....##.
		823 =>	"00111100",	-- ..####..
		824 =>	"00000110",	-- .....##.
		825 =>	"00000110",	-- .....##.
		826 =>	"11000110",	-- ##...##.
		827 =>	"01111100",	-- .#####..
		828 =>	"00000000",	-- ........
		829 =>	"00000000",	-- ........
		830 =>	"00000000",	-- ........
		831 =>	"00000000",	-- ........

		-- char 0x34='4'  
		832 =>	"00000000",	-- ........
		833 =>	"00000000",	-- ........
		834 =>	"00000000",	-- ........
		835 =>	"00001100",	-- ....##..
		836 =>	"00011100",	-- ...###..
		837 =>	"00111100",	-- ..####..
		838 =>	"01101100",	-- .##.##..
		839 =>	"11001100",	-- ##..##..
		840 =>	"11111110",	-- #######.
		841 =>	"00001100",	-- ....##..
		842 =>	"00001100",	-- ....##..
		843 =>	"00011110",	-- ...####.
		844 =>	"00000000",	-- ........
		845 =>	"00000000",	-- ........
		846 =>	"00000000",	-- ........
		847 =>	"00000000",	-- ........

		-- char 0x35='5'  
		848 =>	"00000000",	-- ........
		849 =>	"00000000",	-- ........
		850 =>	"00000000",	-- ........
		851 =>	"11111110",	-- #######.
		852 =>	"11000000",	-- ##......
		853 =>	"11000000",	-- ##......
		854 =>	"11000000",	-- ##......
		855 =>	"11111100",	-- ######..
		856 =>	"00000110",	-- .....##.
		857 =>	"00000110",	-- .....##.
		858 =>	"11000110",	-- ##...##.
		859 =>	"01111100",	-- .#####..
		860 =>	"00000000",	-- ........
		861 =>	"00000000",	-- ........
		862 =>	"00000000",	-- ........
		863 =>	"00000000",	-- ........

		-- char 0x36='6'  
		864 =>	"00000000",	-- ........
		865 =>	"00000000",	-- ........
		866 =>	"00000000",	-- ........
		867 =>	"00111000",	-- ..###...
		868 =>	"01100000",	-- .##.....
		869 =>	"11000000",	-- ##......
		870 =>	"11000000",	-- ##......
		871 =>	"11111100",	-- ######..
		872 =>	"11000110",	-- ##...##.
		873 =>	"11000110",	-- ##...##.
		874 =>	"11000110",	-- ##...##.
		875 =>	"01111100",	-- .#####..
		876 =>	"00000000",	-- ........
		877 =>	"00000000",	-- ........
		878 =>	"00000000",	-- ........
		879 =>	"00000000",	-- ........

		-- char 0x37='7'  
		880 =>	"00000000",	-- ........
		881 =>	"00000000",	-- ........
		882 =>	"00000000",	-- ........
		883 =>	"11111110",	-- #######.
		884 =>	"11000110",	-- ##...##.
		885 =>	"00000110",	-- .....##.
		886 =>	"00001100",	-- ....##..
		887 =>	"00011000",	-- ...##...
		888 =>	"00110000",	-- ..##....
		889 =>	"00110000",	-- ..##....
		890 =>	"00110000",	-- ..##....
		891 =>	"00110000",	-- ..##....
		892 =>	"00000000",	-- ........
		893 =>	"00000000",	-- ........
		894 =>	"00000000",	-- ........
		895 =>	"00000000",	-- ........

		-- char 0x38='8'  
		896 =>	"00000000",	-- ........
		897 =>	"00000000",	-- ........
		898 =>	"00000000",	-- ........
		899 =>	"01111100",	-- .#####..
		900 =>	"11000110",	-- ##...##.
		901 =>	"11000110",	-- ##...##.
		902 =>	"11000110",	-- ##...##.
		903 =>	"01111100",	-- .#####..
		904 =>	"11000110",	-- ##...##.
		905 =>	"11000110",	-- ##...##.
		906 =>	"11000110",	-- ##...##.
		907 =>	"01111100",	-- .#####..
		908 =>	"00000000",	-- ........
		909 =>	"00000000",	-- ........
		910 =>	"00000000",	-- ........
		911 =>	"00000000",	-- ........

		-- char 0x39='9'  
		912 =>	"00000000",	-- ........
		913 =>	"00000000",	-- ........
		914 =>	"00000000",	-- ........
		915 =>	"01111100",	-- .#####..
		916 =>	"11000110",	-- ##...##.
		917 =>	"11000110",	-- ##...##.
		918 =>	"11000110",	-- ##...##.
		919 =>	"01111110",	-- .######.
		920 =>	"00000110",	-- .....##.
		921 =>	"00000110",	-- .....##.
		922 =>	"00001100",	-- ....##..
		923 =>	"01111000",	-- .####...
		924 =>	"00000000",	-- ........
		925 =>	"00000000",	-- ........
		926 =>	"00000000",	-- ........
		927 =>	"00000000",	-- ........

		-- char 0x3a=':'  
		928 =>	"00000000",	-- ........
		929 =>	"00000000",	-- ........
		930 =>	"00000000",	-- ........
		931 =>	"00000000",	-- ........
		932 =>	"00011000",	-- ...##...
		933 =>	"00011000",	-- ...##...
		934 =>	"00000000",	-- ........
		935 =>	"00000000",	-- ........
		936 =>	"00000000",	-- ........
		937 =>	"00011000",	-- ...##...
		938 =>	"00011000",	-- ...##...
		939 =>	"00000000",	-- ........
		940 =>	"00000000",	-- ........
		941 =>	"00000000",	-- ........
		942 =>	"00000000",	-- ........
		943 =>	"00000000",	-- ........

		-- char 0x3b=';'  
		944 =>	"00000000",	-- ........
		945 =>	"00000000",	-- ........
		946 =>	"00000000",	-- ........
		947 =>	"00000000",	-- ........
		948 =>	"00011000",	-- ...##...
		949 =>	"00011000",	-- ...##...
		950 =>	"00000000",	-- ........
		951 =>	"00000000",	-- ........
		952 =>	"00000000",	-- ........
		953 =>	"00011000",	-- ...##...
		954 =>	"00011000",	-- ...##...
		955 =>	"00110000",	-- ..##....
		956 =>	"00000000",	-- ........
		957 =>	"00000000",	-- ........
		958 =>	"00000000",	-- ........
		959 =>	"00000000",	-- ........

		-- char 0x3c='<'  
		960 =>	"00000000",	-- ........
		961 =>	"00000000",	-- ........
		962 =>	"00000000",	-- ........
		963 =>	"00000110",	-- .....##.
		964 =>	"00001100",	-- ....##..
		965 =>	"00011000",	-- ...##...
		966 =>	"00110000",	-- ..##....
		967 =>	"01100000",	-- .##.....
		968 =>	"00110000",	-- ..##....
		969 =>	"00011000",	-- ...##...
		970 =>	"00001100",	-- ....##..
		971 =>	"00000110",	-- .....##.
		972 =>	"00000000",	-- ........
		973 =>	"00000000",	-- ........
		974 =>	"00000000",	-- ........
		975 =>	"00000000",	-- ........

		-- char 0x3d='='  
		976 =>	"00000000",	-- ........
		977 =>	"00000000",	-- ........
		978 =>	"00000000",	-- ........
		979 =>	"00000000",	-- ........
		980 =>	"00000000",	-- ........
		981 =>	"00000000",	-- ........
		982 =>	"01111110",	-- .######.
		983 =>	"00000000",	-- ........
		984 =>	"00000000",	-- ........
		985 =>	"01111110",	-- .######.
		986 =>	"00000000",	-- ........
		987 =>	"00000000",	-- ........
		988 =>	"00000000",	-- ........
		989 =>	"00000000",	-- ........
		990 =>	"00000000",	-- ........
		991 =>	"00000000",	-- ........

		-- char 0x3e='>'  
		992 =>	"00000000",	-- ........
		993 =>	"00000000",	-- ........
		994 =>	"00000000",	-- ........
		995 =>	"01100000",	-- .##.....
		996 =>	"00110000",	-- ..##....
		997 =>	"00011000",	-- ...##...
		998 =>	"00001100",	-- ....##..
		999 =>	"00000110",	-- .....##.
		1000 =>	"00001100",	-- ....##..
		1001 =>	"00011000",	-- ...##...
		1002 =>	"00110000",	-- ..##....
		1003 =>	"01100000",	-- .##.....
		1004 =>	"00000000",	-- ........
		1005 =>	"00000000",	-- ........
		1006 =>	"00000000",	-- ........
		1007 =>	"00000000",	-- ........

		-- char 0x3f='?'  
		1008 =>	"00000000",	-- ........
		1009 =>	"00000000",	-- ........
		1010 =>	"00000000",	-- ........
		1011 =>	"01111100",	-- .#####..
		1012 =>	"11000110",	-- ##...##.
		1013 =>	"11000110",	-- ##...##.
		1014 =>	"00001100",	-- ....##..
		1015 =>	"00011000",	-- ...##...
		1016 =>	"00011000",	-- ...##...
		1017 =>	"00000000",	-- ........
		1018 =>	"00011000",	-- ...##...
		1019 =>	"00011000",	-- ...##...
		1020 =>	"00000000",	-- ........
		1021 =>	"00000000",	-- ........
		1022 =>	"00000000",	-- ........
		1023 =>	"00000000",	-- ........

		-- char 0x40='@'  
		1024 =>	"00000000",	-- ........
		1025 =>	"00000000",	-- ........
		1026 =>	"00000000",	-- ........
		1027 =>	"01111100",	-- .#####..
		1028 =>	"11000110",	-- ##...##.
		1029 =>	"11000110",	-- ##...##.
		1030 =>	"11011110",	-- ##.####.
		1031 =>	"11011110",	-- ##.####.
		1032 =>	"11011110",	-- ##.####.
		1033 =>	"11011100",	-- ##.###..
		1034 =>	"11000000",	-- ##......
		1035 =>	"01111100",	-- .#####..
		1036 =>	"00000000",	-- ........
		1037 =>	"00000000",	-- ........
		1038 =>	"00000000",	-- ........
		1039 =>	"00000000",	-- ........

		-- char 0x41='A'  
		1040 =>	"00000000",	-- ........
		1041 =>	"00000000",	-- ........
		1042 =>	"00000000",	-- ........
		1043 =>	"00010000",	-- ...#....
		1044 =>	"00111000",	-- ..###...
		1045 =>	"01101100",	-- .##.##..
		1046 =>	"11000110",	-- ##...##.
		1047 =>	"11000110",	-- ##...##.
		1048 =>	"11111110",	-- #######.
		1049 =>	"11000110",	-- ##...##.
		1050 =>	"11000110",	-- ##...##.
		1051 =>	"11000110",	-- ##...##.
		1052 =>	"00000000",	-- ........
		1053 =>	"00000000",	-- ........
		1054 =>	"00000000",	-- ........
		1055 =>	"00000000",	-- ........

		-- char 0x42='B'  
		1056 =>	"00000000",	-- ........
		1057 =>	"00000000",	-- ........
		1058 =>	"00000000",	-- ........
		1059 =>	"11111100",	-- ######..
		1060 =>	"01100110",	-- .##..##.
		1061 =>	"01100110",	-- .##..##.
		1062 =>	"01100110",	-- .##..##.
		1063 =>	"01111100",	-- .#####..
		1064 =>	"01100110",	-- .##..##.
		1065 =>	"01100110",	-- .##..##.
		1066 =>	"01100110",	-- .##..##.
		1067 =>	"11111100",	-- ######..
		1068 =>	"00000000",	-- ........
		1069 =>	"00000000",	-- ........
		1070 =>	"00000000",	-- ........
		1071 =>	"00000000",	-- ........

		-- char 0x43='C'  
		1072 =>	"00000000",	-- ........
		1073 =>	"00000000",	-- ........
		1074 =>	"00000000",	-- ........
		1075 =>	"00111100",	-- ..####..
		1076 =>	"01100110",	-- .##..##.
		1077 =>	"11000010",	-- ##....#.
		1078 =>	"11000000",	-- ##......
		1079 =>	"11000000",	-- ##......
		1080 =>	"11000000",	-- ##......
		1081 =>	"11000010",	-- ##....#.
		1082 =>	"01100110",	-- .##..##.
		1083 =>	"00111100",	-- ..####..
		1084 =>	"00000000",	-- ........
		1085 =>	"00000000",	-- ........
		1086 =>	"00000000",	-- ........
		1087 =>	"00000000",	-- ........

		-- char 0x44='D'  
		1088 =>	"00000000",	-- ........
		1089 =>	"00000000",	-- ........
		1090 =>	"00000000",	-- ........
		1091 =>	"11111000",	-- #####...
		1092 =>	"01101100",	-- .##.##..
		1093 =>	"01100110",	-- .##..##.
		1094 =>	"01100110",	-- .##..##.
		1095 =>	"01100110",	-- .##..##.
		1096 =>	"01100110",	-- .##..##.
		1097 =>	"01100110",	-- .##..##.
		1098 =>	"01101100",	-- .##.##..
		1099 =>	"11111000",	-- #####...
		1100 =>	"00000000",	-- ........
		1101 =>	"00000000",	-- ........
		1102 =>	"00000000",	-- ........
		1103 =>	"00000000",	-- ........

		-- char 0x45='E'  
		1104 =>	"00000000",	-- ........
		1105 =>	"00000000",	-- ........
		1106 =>	"00000000",	-- ........
		1107 =>	"11111110",	-- #######.
		1108 =>	"01100110",	-- .##..##.
		1109 =>	"01100010",	-- .##...#.
		1110 =>	"01101000",	-- .##.#...
		1111 =>	"01111000",	-- .####...
		1112 =>	"01101000",	-- .##.#...
		1113 =>	"01100010",	-- .##...#.
		1114 =>	"01100110",	-- .##..##.
		1115 =>	"11111110",	-- #######.
		1116 =>	"00000000",	-- ........
		1117 =>	"00000000",	-- ........
		1118 =>	"00000000",	-- ........
		1119 =>	"00000000",	-- ........

		-- char 0x46='F'  
		1120 =>	"00000000",	-- ........
		1121 =>	"00000000",	-- ........
		1122 =>	"00000000",	-- ........
		1123 =>	"11111110",	-- #######.
		1124 =>	"01100110",	-- .##..##.
		1125 =>	"01100010",	-- .##...#.
		1126 =>	"01101000",	-- .##.#...
		1127 =>	"01111000",	-- .####...
		1128 =>	"01101000",	-- .##.#...
		1129 =>	"01100000",	-- .##.....
		1130 =>	"01100000",	-- .##.....
		1131 =>	"11110000",	-- ####....
		1132 =>	"00000000",	-- ........
		1133 =>	"00000000",	-- ........
		1134 =>	"00000000",	-- ........
		1135 =>	"00000000",	-- ........

		-- char 0x47='G'  
		1136 =>	"00000000",	-- ........
		1137 =>	"00000000",	-- ........
		1138 =>	"00000000",	-- ........
		1139 =>	"00111100",	-- ..####..
		1140 =>	"01100110",	-- .##..##.
		1141 =>	"11000010",	-- ##....#.
		1142 =>	"11000000",	-- ##......
		1143 =>	"11000000",	-- ##......
		1144 =>	"11011110",	-- ##.####.
		1145 =>	"11000110",	-- ##...##.
		1146 =>	"01100110",	-- .##..##.
		1147 =>	"00111010",	-- ..###.#.
		1148 =>	"00000000",	-- ........
		1149 =>	"00000000",	-- ........
		1150 =>	"00000000",	-- ........
		1151 =>	"00000000",	-- ........

		-- char 0x48='H'  
		1152 =>	"00000000",	-- ........
		1153 =>	"00000000",	-- ........
		1154 =>	"00000000",	-- ........
		1155 =>	"11000110",	-- ##...##.
		1156 =>	"11000110",	-- ##...##.
		1157 =>	"11000110",	-- ##...##.
		1158 =>	"11000110",	-- ##...##.
		1159 =>	"11111110",	-- #######.
		1160 =>	"11000110",	-- ##...##.
		1161 =>	"11000110",	-- ##...##.
		1162 =>	"11000110",	-- ##...##.
		1163 =>	"11000110",	-- ##...##.
		1164 =>	"00000000",	-- ........
		1165 =>	"00000000",	-- ........
		1166 =>	"00000000",	-- ........
		1167 =>	"00000000",	-- ........

		-- char 0x49='I'  
		1168 =>	"00000000",	-- ........
		1169 =>	"00000000",	-- ........
		1170 =>	"00000000",	-- ........
		1171 =>	"00111100",	-- ..####..
		1172 =>	"00011000",	-- ...##...
		1173 =>	"00011000",	-- ...##...
		1174 =>	"00011000",	-- ...##...
		1175 =>	"00011000",	-- ...##...
		1176 =>	"00011000",	-- ...##...
		1177 =>	"00011000",	-- ...##...
		1178 =>	"00011000",	-- ...##...
		1179 =>	"00111100",	-- ..####..
		1180 =>	"00000000",	-- ........
		1181 =>	"00000000",	-- ........
		1182 =>	"00000000",	-- ........
		1183 =>	"00000000",	-- ........

		-- char 0x4a='J'  
		1184 =>	"00000000",	-- ........
		1185 =>	"00000000",	-- ........
		1186 =>	"00000000",	-- ........
		1187 =>	"00011110",	-- ...####.
		1188 =>	"00001100",	-- ....##..
		1189 =>	"00001100",	-- ....##..
		1190 =>	"00001100",	-- ....##..
		1191 =>	"00001100",	-- ....##..
		1192 =>	"00001100",	-- ....##..
		1193 =>	"11001100",	-- ##..##..
		1194 =>	"11001100",	-- ##..##..
		1195 =>	"01111000",	-- .####...
		1196 =>	"00000000",	-- ........
		1197 =>	"00000000",	-- ........
		1198 =>	"00000000",	-- ........
		1199 =>	"00000000",	-- ........

		-- char 0x4b='K'  
		1200 =>	"00000000",	-- ........
		1201 =>	"00000000",	-- ........
		1202 =>	"00000000",	-- ........
		1203 =>	"11100110",	-- ###..##.
		1204 =>	"01100110",	-- .##..##.
		1205 =>	"01101100",	-- .##.##..
		1206 =>	"01101100",	-- .##.##..
		1207 =>	"01111000",	-- .####...
		1208 =>	"01101100",	-- .##.##..
		1209 =>	"01101100",	-- .##.##..
		1210 =>	"01100110",	-- .##..##.
		1211 =>	"11100110",	-- ###..##.
		1212 =>	"00000000",	-- ........
		1213 =>	"00000000",	-- ........
		1214 =>	"00000000",	-- ........
		1215 =>	"00000000",	-- ........

		-- char 0x4c='L'  
		1216 =>	"00000000",	-- ........
		1217 =>	"00000000",	-- ........
		1218 =>	"00000000",	-- ........
		1219 =>	"11110000",	-- ####....
		1220 =>	"01100000",	-- .##.....
		1221 =>	"01100000",	-- .##.....
		1222 =>	"01100000",	-- .##.....
		1223 =>	"01100000",	-- .##.....
		1224 =>	"01100000",	-- .##.....
		1225 =>	"01100010",	-- .##...#.
		1226 =>	"01100110",	-- .##..##.
		1227 =>	"11111110",	-- #######.
		1228 =>	"00000000",	-- ........
		1229 =>	"00000000",	-- ........
		1230 =>	"00000000",	-- ........
		1231 =>	"00000000",	-- ........

		-- char 0x4d='M'  
		1232 =>	"00000000",	-- ........
		1233 =>	"00000000",	-- ........
		1234 =>	"00000000",	-- ........
		1235 =>	"11000110",	-- ##...##.
		1236 =>	"11101110",	-- ###.###.
		1237 =>	"11111110",	-- #######.
		1238 =>	"11111110",	-- #######.
		1239 =>	"11010110",	-- ##.#.##.
		1240 =>	"11000110",	-- ##...##.
		1241 =>	"11000110",	-- ##...##.
		1242 =>	"11000110",	-- ##...##.
		1243 =>	"11000110",	-- ##...##.
		1244 =>	"00000000",	-- ........
		1245 =>	"00000000",	-- ........
		1246 =>	"00000000",	-- ........
		1247 =>	"00000000",	-- ........

		-- char 0x4e='N'  
		1248 =>	"00000000",	-- ........
		1249 =>	"00000000",	-- ........
		1250 =>	"00000000",	-- ........
		1251 =>	"11000110",	-- ##...##.
		1252 =>	"11100110",	-- ###..##.
		1253 =>	"11110110",	-- ####.##.
		1254 =>	"11111110",	-- #######.
		1255 =>	"11011110",	-- ##.####.
		1256 =>	"11001110",	-- ##..###.
		1257 =>	"11000110",	-- ##...##.
		1258 =>	"11000110",	-- ##...##.
		1259 =>	"11000110",	-- ##...##.
		1260 =>	"00000000",	-- ........
		1261 =>	"00000000",	-- ........
		1262 =>	"00000000",	-- ........
		1263 =>	"00000000",	-- ........

		-- char 0x4f='O'  
		1264 =>	"00000000",	-- ........
		1265 =>	"00000000",	-- ........
		1266 =>	"00000000",	-- ........
		1267 =>	"00111000",	-- ..###...
		1268 =>	"01101100",	-- .##.##..
		1269 =>	"11000110",	-- ##...##.
		1270 =>	"11000110",	-- ##...##.
		1271 =>	"11000110",	-- ##...##.
		1272 =>	"11000110",	-- ##...##.
		1273 =>	"11000110",	-- ##...##.
		1274 =>	"01101100",	-- .##.##..
		1275 =>	"00111000",	-- ..###...
		1276 =>	"00000000",	-- ........
		1277 =>	"00000000",	-- ........
		1278 =>	"00000000",	-- ........
		1279 =>	"00000000",	-- ........

		-- char 0x50='P'  
		1280 =>	"00000000",	-- ........
		1281 =>	"00000000",	-- ........
		1282 =>	"00000000",	-- ........
		1283 =>	"11111100",	-- ######..
		1284 =>	"01100110",	-- .##..##.
		1285 =>	"01100110",	-- .##..##.
		1286 =>	"01100110",	-- .##..##.
		1287 =>	"01111100",	-- .#####..
		1288 =>	"01100000",	-- .##.....
		1289 =>	"01100000",	-- .##.....
		1290 =>	"01100000",	-- .##.....
		1291 =>	"11110000",	-- ####....
		1292 =>	"00000000",	-- ........
		1293 =>	"00000000",	-- ........
		1294 =>	"00000000",	-- ........
		1295 =>	"00000000",	-- ........

		-- char 0x51='Q'  
		1296 =>	"00000000",	-- ........
		1297 =>	"00000000",	-- ........
		1298 =>	"00000000",	-- ........
		1299 =>	"01111100",	-- .#####..
		1300 =>	"11000110",	-- ##...##.
		1301 =>	"11000110",	-- ##...##.
		1302 =>	"11000110",	-- ##...##.
		1303 =>	"11000110",	-- ##...##.
		1304 =>	"11010110",	-- ##.#.##.
		1305 =>	"11011110",	-- ##.####.
		1306 =>	"01111100",	-- .#####..
		1307 =>	"00001100",	-- ....##..
		1308 =>	"00001110",	-- ....###.
		1309 =>	"00000000",	-- ........
		1310 =>	"00000000",	-- ........
		1311 =>	"00000000",	-- ........

		-- char 0x52='R'  
		1312 =>	"00000000",	-- ........
		1313 =>	"00000000",	-- ........
		1314 =>	"00000000",	-- ........
		1315 =>	"11111100",	-- ######..
		1316 =>	"01100110",	-- .##..##.
		1317 =>	"01100110",	-- .##..##.
		1318 =>	"01100110",	-- .##..##.
		1319 =>	"01111100",	-- .#####..
		1320 =>	"01101100",	-- .##.##..
		1321 =>	"01100110",	-- .##..##.
		1322 =>	"01100110",	-- .##..##.
		1323 =>	"11100110",	-- ###..##.
		1324 =>	"00000000",	-- ........
		1325 =>	"00000000",	-- ........
		1326 =>	"00000000",	-- ........
		1327 =>	"00000000",	-- ........

		-- char 0x53='S'  
		1328 =>	"00000000",	-- ........
		1329 =>	"00000000",	-- ........
		1330 =>	"00000000",	-- ........
		1331 =>	"01111100",	-- .#####..
		1332 =>	"11000110",	-- ##...##.
		1333 =>	"11000110",	-- ##...##.
		1334 =>	"01100000",	-- .##.....
		1335 =>	"00111000",	-- ..###...
		1336 =>	"00001100",	-- ....##..
		1337 =>	"11000110",	-- ##...##.
		1338 =>	"11000110",	-- ##...##.
		1339 =>	"01111100",	-- .#####..
		1340 =>	"00000000",	-- ........
		1341 =>	"00000000",	-- ........
		1342 =>	"00000000",	-- ........
		1343 =>	"00000000",	-- ........

		-- char 0x54='T'  
		1344 =>	"00000000",	-- ........
		1345 =>	"00000000",	-- ........
		1346 =>	"00000000",	-- ........
		1347 =>	"01111110",	-- .######.
		1348 =>	"01111110",	-- .######.
		1349 =>	"01011010",	-- .#.##.#.
		1350 =>	"00011000",	-- ...##...
		1351 =>	"00011000",	-- ...##...
		1352 =>	"00011000",	-- ...##...
		1353 =>	"00011000",	-- ...##...
		1354 =>	"00011000",	-- ...##...
		1355 =>	"00111100",	-- ..####..
		1356 =>	"00000000",	-- ........
		1357 =>	"00000000",	-- ........
		1358 =>	"00000000",	-- ........
		1359 =>	"00000000",	-- ........

		-- char 0x55='U'  
		1360 =>	"00000000",	-- ........
		1361 =>	"00000000",	-- ........
		1362 =>	"00000000",	-- ........
		1363 =>	"11000110",	-- ##...##.
		1364 =>	"11000110",	-- ##...##.
		1365 =>	"11000110",	-- ##...##.
		1366 =>	"11000110",	-- ##...##.
		1367 =>	"11000110",	-- ##...##.
		1368 =>	"11000110",	-- ##...##.
		1369 =>	"11000110",	-- ##...##.
		1370 =>	"11000110",	-- ##...##.
		1371 =>	"01111100",	-- .#####..
		1372 =>	"00000000",	-- ........
		1373 =>	"00000000",	-- ........
		1374 =>	"00000000",	-- ........
		1375 =>	"00000000",	-- ........

		-- char 0x56='V'  
		1376 =>	"00000000",	-- ........
		1377 =>	"00000000",	-- ........
		1378 =>	"00000000",	-- ........
		1379 =>	"11000110",	-- ##...##.
		1380 =>	"11000110",	-- ##...##.
		1381 =>	"11000110",	-- ##...##.
		1382 =>	"11000110",	-- ##...##.
		1383 =>	"11000110",	-- ##...##.
		1384 =>	"11000110",	-- ##...##.
		1385 =>	"01101100",	-- .##.##..
		1386 =>	"00111000",	-- ..###...
		1387 =>	"00010000",	-- ...#....
		1388 =>	"00000000",	-- ........
		1389 =>	"00000000",	-- ........
		1390 =>	"00000000",	-- ........
		1391 =>	"00000000",	-- ........

		-- char 0x57='W'  
		1392 =>	"00000000",	-- ........
		1393 =>	"00000000",	-- ........
		1394 =>	"00000000",	-- ........
		1395 =>	"11000110",	-- ##...##.
		1396 =>	"11000110",	-- ##...##.
		1397 =>	"11000110",	-- ##...##.
		1398 =>	"11000110",	-- ##...##.
		1399 =>	"11010110",	-- ##.#.##.
		1400 =>	"11010110",	-- ##.#.##.
		1401 =>	"11111110",	-- #######.
		1402 =>	"01111100",	-- .#####..
		1403 =>	"01101100",	-- .##.##..
		1404 =>	"00000000",	-- ........
		1405 =>	"00000000",	-- ........
		1406 =>	"00000000",	-- ........
		1407 =>	"00000000",	-- ........

		-- char 0x58='X'  
		1408 =>	"00000000",	-- ........
		1409 =>	"00000000",	-- ........
		1410 =>	"00000000",	-- ........
		1411 =>	"11000110",	-- ##...##.
		1412 =>	"11000110",	-- ##...##.
		1413 =>	"01101100",	-- .##.##..
		1414 =>	"00111000",	-- ..###...
		1415 =>	"00111000",	-- ..###...
		1416 =>	"00111000",	-- ..###...
		1417 =>	"01101100",	-- .##.##..
		1418 =>	"11000110",	-- ##...##.
		1419 =>	"11000110",	-- ##...##.
		1420 =>	"00000000",	-- ........
		1421 =>	"00000000",	-- ........
		1422 =>	"00000000",	-- ........
		1423 =>	"00000000",	-- ........

		-- char 0x59='Y'  
		1424 =>	"00000000",	-- ........
		1425 =>	"00000000",	-- ........
		1426 =>	"00000000",	-- ........
		1427 =>	"01100110",	-- .##..##.
		1428 =>	"01100110",	-- .##..##.
		1429 =>	"01100110",	-- .##..##.
		1430 =>	"01100110",	-- .##..##.
		1431 =>	"00111100",	-- ..####..
		1432 =>	"00011000",	-- ...##...
		1433 =>	"00011000",	-- ...##...
		1434 =>	"00011000",	-- ...##...
		1435 =>	"00111100",	-- ..####..
		1436 =>	"00000000",	-- ........
		1437 =>	"00000000",	-- ........
		1438 =>	"00000000",	-- ........
		1439 =>	"00000000",	-- ........

		-- char 0x5a='Z'  
		1440 =>	"00000000",	-- ........
		1441 =>	"00000000",	-- ........
		1442 =>	"00000000",	-- ........
		1443 =>	"11111110",	-- #######.
		1444 =>	"11000110",	-- ##...##.
		1445 =>	"10001100",	-- #...##..
		1446 =>	"00011000",	-- ...##...
		1447 =>	"00110000",	-- ..##....
		1448 =>	"01100000",	-- .##.....
		1449 =>	"11000010",	-- ##....#.
		1450 =>	"11000110",	-- ##...##.
		1451 =>	"11111110",	-- #######.
		1452 =>	"00000000",	-- ........
		1453 =>	"00000000",	-- ........
		1454 =>	"00000000",	-- ........
		1455 =>	"00000000",	-- ........

		-- char 0x5b='['  
		1456 =>	"00000000",	-- ........
		1457 =>	"00000000",	-- ........
		1458 =>	"00000000",	-- ........
		1459 =>	"00111100",	-- ..####..
		1460 =>	"00110000",	-- ..##....
		1461 =>	"00110000",	-- ..##....
		1462 =>	"00110000",	-- ..##....
		1463 =>	"00110000",	-- ..##....
		1464 =>	"00110000",	-- ..##....
		1465 =>	"00110000",	-- ..##....
		1466 =>	"00110000",	-- ..##....
		1467 =>	"00111100",	-- ..####..
		1468 =>	"00000000",	-- ........
		1469 =>	"00000000",	-- ........
		1470 =>	"00000000",	-- ........
		1471 =>	"00000000",	-- ........

		-- char 0x5c='\\' 
		1472 =>	"00000000",	-- ........
		1473 =>	"00000000",	-- ........
		1474 =>	"00000000",	-- ........
		1475 =>	"10000000",	-- #.......
		1476 =>	"11000000",	-- ##......
		1477 =>	"11100000",	-- ###.....
		1478 =>	"01110000",	-- .###....
		1479 =>	"00111000",	-- ..###...
		1480 =>	"00011100",	-- ...###..
		1481 =>	"00001110",	-- ....###.
		1482 =>	"00000110",	-- .....##.
		1483 =>	"00000010",	-- ......#.
		1484 =>	"00000000",	-- ........
		1485 =>	"00000000",	-- ........
		1486 =>	"00000000",	-- ........
		1487 =>	"00000000",	-- ........

		-- char 0x5d=']'  
		1488 =>	"00000000",	-- ........
		1489 =>	"00000000",	-- ........
		1490 =>	"00000000",	-- ........
		1491 =>	"00111100",	-- ..####..
		1492 =>	"00001100",	-- ....##..
		1493 =>	"00001100",	-- ....##..
		1494 =>	"00001100",	-- ....##..
		1495 =>	"00001100",	-- ....##..
		1496 =>	"00001100",	-- ....##..
		1497 =>	"00001100",	-- ....##..
		1498 =>	"00001100",	-- ....##..
		1499 =>	"00111100",	-- ..####..
		1500 =>	"00000000",	-- ........
		1501 =>	"00000000",	-- ........
		1502 =>	"00000000",	-- ........
		1503 =>	"00000000",	-- ........

		-- char 0x5e='^'  
		1504 =>	"00000000",	-- ........
		1505 =>	"00010000",	-- ...#....
		1506 =>	"00111000",	-- ..###...
		1507 =>	"01101100",	-- .##.##..
		1508 =>	"11000110",	-- ##...##.
		1509 =>	"00000000",	-- ........
		1510 =>	"00000000",	-- ........
		1511 =>	"00000000",	-- ........
		1512 =>	"00000000",	-- ........
		1513 =>	"00000000",	-- ........
		1514 =>	"00000000",	-- ........
		1515 =>	"00000000",	-- ........
		1516 =>	"00000000",	-- ........
		1517 =>	"00000000",	-- ........
		1518 =>	"00000000",	-- ........
		1519 =>	"00000000",	-- ........

		-- char 0x5f='_'  
		1520 =>	"00000000",	-- ........
		1521 =>	"00000000",	-- ........
		1522 =>	"00000000",	-- ........
		1523 =>	"00000000",	-- ........
		1524 =>	"00000000",	-- ........
		1525 =>	"00000000",	-- ........
		1526 =>	"00000000",	-- ........
		1527 =>	"00000000",	-- ........
		1528 =>	"00000000",	-- ........
		1529 =>	"00000000",	-- ........
		1530 =>	"00000000",	-- ........
		1531 =>	"00000000",	-- ........
		1532 =>	"00000000",	-- ........
		1533 =>	"11111111",	-- ########
		1534 =>	"00000000",	-- ........
		1535 =>	"00000000",	-- ........

		-- char 0x60='`'  
		1536 =>	"00000000",	-- ........
		1537 =>	"00110000",	-- ..##....
		1538 =>	"00110000",	-- ..##....
		1539 =>	"00011000",	-- ...##...
		1540 =>	"00000000",	-- ........
		1541 =>	"00000000",	-- ........
		1542 =>	"00000000",	-- ........
		1543 =>	"00000000",	-- ........
		1544 =>	"00000000",	-- ........
		1545 =>	"00000000",	-- ........
		1546 =>	"00000000",	-- ........
		1547 =>	"00000000",	-- ........
		1548 =>	"00000000",	-- ........
		1549 =>	"00000000",	-- ........
		1550 =>	"00000000",	-- ........
		1551 =>	"00000000",	-- ........

		-- char 0x61='a'  
		1552 =>	"00000000",	-- ........
		1553 =>	"00000000",	-- ........
		1554 =>	"00000000",	-- ........
		1555 =>	"00000000",	-- ........
		1556 =>	"00000000",	-- ........
		1557 =>	"00000000",	-- ........
		1558 =>	"01111000",	-- .####...
		1559 =>	"00001100",	-- ....##..
		1560 =>	"01111100",	-- .#####..
		1561 =>	"11001100",	-- ##..##..
		1562 =>	"11001100",	-- ##..##..
		1563 =>	"01110110",	-- .###.##.
		1564 =>	"00000000",	-- ........
		1565 =>	"00000000",	-- ........
		1566 =>	"00000000",	-- ........
		1567 =>	"00000000",	-- ........

		-- char 0x62='b'  
		1568 =>	"00000000",	-- ........
		1569 =>	"00000000",	-- ........
		1570 =>	"00000000",	-- ........
		1571 =>	"11100000",	-- ###.....
		1572 =>	"01100000",	-- .##.....
		1573 =>	"01100000",	-- .##.....
		1574 =>	"01111000",	-- .####...
		1575 =>	"01101100",	-- .##.##..
		1576 =>	"01100110",	-- .##..##.
		1577 =>	"01100110",	-- .##..##.
		1578 =>	"01100110",	-- .##..##.
		1579 =>	"01111100",	-- .#####..
		1580 =>	"00000000",	-- ........
		1581 =>	"00000000",	-- ........
		1582 =>	"00000000",	-- ........
		1583 =>	"00000000",	-- ........

		-- char 0x63='c'  
		1584 =>	"00000000",	-- ........
		1585 =>	"00000000",	-- ........
		1586 =>	"00000000",	-- ........
		1587 =>	"00000000",	-- ........
		1588 =>	"00000000",	-- ........
		1589 =>	"00000000",	-- ........
		1590 =>	"01111100",	-- .#####..
		1591 =>	"11000110",	-- ##...##.
		1592 =>	"11000000",	-- ##......
		1593 =>	"11000000",	-- ##......
		1594 =>	"11000110",	-- ##...##.
		1595 =>	"01111100",	-- .#####..
		1596 =>	"00000000",	-- ........
		1597 =>	"00000000",	-- ........
		1598 =>	"00000000",	-- ........
		1599 =>	"00000000",	-- ........

		-- char 0x64='d'  
		1600 =>	"00000000",	-- ........
		1601 =>	"00000000",	-- ........
		1602 =>	"00000000",	-- ........
		1603 =>	"00011100",	-- ...###..
		1604 =>	"00001100",	-- ....##..
		1605 =>	"00001100",	-- ....##..
		1606 =>	"00111100",	-- ..####..
		1607 =>	"01101100",	-- .##.##..
		1608 =>	"11001100",	-- ##..##..
		1609 =>	"11001100",	-- ##..##..
		1610 =>	"11001100",	-- ##..##..
		1611 =>	"01110110",	-- .###.##.
		1612 =>	"00000000",	-- ........
		1613 =>	"00000000",	-- ........
		1614 =>	"00000000",	-- ........
		1615 =>	"00000000",	-- ........

		-- char 0x65='e'  
		1616 =>	"00000000",	-- ........
		1617 =>	"00000000",	-- ........
		1618 =>	"00000000",	-- ........
		1619 =>	"00000000",	-- ........
		1620 =>	"00000000",	-- ........
		1621 =>	"00000000",	-- ........
		1622 =>	"01111100",	-- .#####..
		1623 =>	"11000110",	-- ##...##.
		1624 =>	"11111110",	-- #######.
		1625 =>	"11000000",	-- ##......
		1626 =>	"11000110",	-- ##...##.
		1627 =>	"01111100",	-- .#####..
		1628 =>	"00000000",	-- ........
		1629 =>	"00000000",	-- ........
		1630 =>	"00000000",	-- ........
		1631 =>	"00000000",	-- ........

		-- char 0x66='f'  
		1632 =>	"00000000",	-- ........
		1633 =>	"00000000",	-- ........
		1634 =>	"00000000",	-- ........
		1635 =>	"00111000",	-- ..###...
		1636 =>	"01101100",	-- .##.##..
		1637 =>	"01100100",	-- .##..#..
		1638 =>	"01100000",	-- .##.....
		1639 =>	"11110000",	-- ####....
		1640 =>	"01100000",	-- .##.....
		1641 =>	"01100000",	-- .##.....
		1642 =>	"01100000",	-- .##.....
		1643 =>	"11110000",	-- ####....
		1644 =>	"00000000",	-- ........
		1645 =>	"00000000",	-- ........
		1646 =>	"00000000",	-- ........
		1647 =>	"00000000",	-- ........

		-- char 0x67='g'  
		1648 =>	"00000000",	-- ........
		1649 =>	"00000000",	-- ........
		1650 =>	"00000000",	-- ........
		1651 =>	"00000000",	-- ........
		1652 =>	"00000000",	-- ........
		1653 =>	"00000000",	-- ........
		1654 =>	"01110110",	-- .###.##.
		1655 =>	"11001100",	-- ##..##..
		1656 =>	"11001100",	-- ##..##..
		1657 =>	"11001100",	-- ##..##..
		1658 =>	"01111100",	-- .#####..
		1659 =>	"00001100",	-- ....##..
		1660 =>	"11001100",	-- ##..##..
		1661 =>	"01111000",	-- .####...
		1662 =>	"00000000",	-- ........
		1663 =>	"00000000",	-- ........

		-- char 0x68='h'  
		1664 =>	"00000000",	-- ........
		1665 =>	"00000000",	-- ........
		1666 =>	"00000000",	-- ........
		1667 =>	"11100000",	-- ###.....
		1668 =>	"01100000",	-- .##.....
		1669 =>	"01100000",	-- .##.....
		1670 =>	"01101100",	-- .##.##..
		1671 =>	"01110110",	-- .###.##.
		1672 =>	"01100110",	-- .##..##.
		1673 =>	"01100110",	-- .##..##.
		1674 =>	"01100110",	-- .##..##.
		1675 =>	"11100110",	-- ###..##.
		1676 =>	"00000000",	-- ........
		1677 =>	"00000000",	-- ........
		1678 =>	"00000000",	-- ........
		1679 =>	"00000000",	-- ........

		-- char 0x69='i'  
		1680 =>	"00000000",	-- ........
		1681 =>	"00000000",	-- ........
		1682 =>	"00000000",	-- ........
		1683 =>	"00011000",	-- ...##...
		1684 =>	"00011000",	-- ...##...
		1685 =>	"00000000",	-- ........
		1686 =>	"00111000",	-- ..###...
		1687 =>	"00011000",	-- ...##...
		1688 =>	"00011000",	-- ...##...
		1689 =>	"00011000",	-- ...##...
		1690 =>	"00011000",	-- ...##...
		1691 =>	"00111100",	-- ..####..
		1692 =>	"00000000",	-- ........
		1693 =>	"00000000",	-- ........
		1694 =>	"00000000",	-- ........
		1695 =>	"00000000",	-- ........

		-- char 0x6a='j'  
		1696 =>	"00000000",	-- ........
		1697 =>	"00000000",	-- ........
		1698 =>	"00000000",	-- ........
		1699 =>	"00000110",	-- .....##.
		1700 =>	"00000110",	-- .....##.
		1701 =>	"00000000",	-- ........
		1702 =>	"00001110",	-- ....###.
		1703 =>	"00000110",	-- .....##.
		1704 =>	"00000110",	-- .....##.
		1705 =>	"00000110",	-- .....##.
		1706 =>	"00000110",	-- .....##.
		1707 =>	"01100110",	-- .##..##.
		1708 =>	"01100110",	-- .##..##.
		1709 =>	"00111100",	-- ..####..
		1710 =>	"00000000",	-- ........
		1711 =>	"00000000",	-- ........

		-- char 0x6b='k'  
		1712 =>	"00000000",	-- ........
		1713 =>	"00000000",	-- ........
		1714 =>	"00000000",	-- ........
		1715 =>	"11100000",	-- ###.....
		1716 =>	"01100000",	-- .##.....
		1717 =>	"01100000",	-- .##.....
		1718 =>	"01100110",	-- .##..##.
		1719 =>	"01101100",	-- .##.##..
		1720 =>	"01111000",	-- .####...
		1721 =>	"01101100",	-- .##.##..
		1722 =>	"01100110",	-- .##..##.
		1723 =>	"11100110",	-- ###..##.
		1724 =>	"00000000",	-- ........
		1725 =>	"00000000",	-- ........
		1726 =>	"00000000",	-- ........
		1727 =>	"00000000",	-- ........

		-- char 0x6c='l'  
		1728 =>	"00000000",	-- ........
		1729 =>	"00000000",	-- ........
		1730 =>	"00000000",	-- ........
		1731 =>	"00111000",	-- ..###...
		1732 =>	"00011000",	-- ...##...
		1733 =>	"00011000",	-- ...##...
		1734 =>	"00011000",	-- ...##...
		1735 =>	"00011000",	-- ...##...
		1736 =>	"00011000",	-- ...##...
		1737 =>	"00011000",	-- ...##...
		1738 =>	"00011000",	-- ...##...
		1739 =>	"00111100",	-- ..####..
		1740 =>	"00000000",	-- ........
		1741 =>	"00000000",	-- ........
		1742 =>	"00000000",	-- ........
		1743 =>	"00000000",	-- ........

		-- char 0x6d='m'  
		1744 =>	"00000000",	-- ........
		1745 =>	"00000000",	-- ........
		1746 =>	"00000000",	-- ........
		1747 =>	"00000000",	-- ........
		1748 =>	"00000000",	-- ........
		1749 =>	"00000000",	-- ........
		1750 =>	"11101100",	-- ###.##..
		1751 =>	"11111110",	-- #######.
		1752 =>	"11010110",	-- ##.#.##.
		1753 =>	"11010110",	-- ##.#.##.
		1754 =>	"11010110",	-- ##.#.##.
		1755 =>	"11000110",	-- ##...##.
		1756 =>	"00000000",	-- ........
		1757 =>	"00000000",	-- ........
		1758 =>	"00000000",	-- ........
		1759 =>	"00000000",	-- ........

		-- char 0x6e='n'  
		1760 =>	"00000000",	-- ........
		1761 =>	"00000000",	-- ........
		1762 =>	"00000000",	-- ........
		1763 =>	"00000000",	-- ........
		1764 =>	"00000000",	-- ........
		1765 =>	"00000000",	-- ........
		1766 =>	"11011100",	-- ##.###..
		1767 =>	"01100110",	-- .##..##.
		1768 =>	"01100110",	-- .##..##.
		1769 =>	"01100110",	-- .##..##.
		1770 =>	"01100110",	-- .##..##.
		1771 =>	"01100110",	-- .##..##.
		1772 =>	"00000000",	-- ........
		1773 =>	"00000000",	-- ........
		1774 =>	"00000000",	-- ........
		1775 =>	"00000000",	-- ........

		-- char 0x6f='o'  
		1776 =>	"00000000",	-- ........
		1777 =>	"00000000",	-- ........
		1778 =>	"00000000",	-- ........
		1779 =>	"00000000",	-- ........
		1780 =>	"00000000",	-- ........
		1781 =>	"00000000",	-- ........
		1782 =>	"01111100",	-- .#####..
		1783 =>	"11000110",	-- ##...##.
		1784 =>	"11000110",	-- ##...##.
		1785 =>	"11000110",	-- ##...##.
		1786 =>	"11000110",	-- ##...##.
		1787 =>	"01111100",	-- .#####..
		1788 =>	"00000000",	-- ........
		1789 =>	"00000000",	-- ........
		1790 =>	"00000000",	-- ........
		1791 =>	"00000000",	-- ........

		-- char 0x70='p'  
		1792 =>	"00000000",	-- ........
		1793 =>	"00000000",	-- ........
		1794 =>	"00000000",	-- ........
		1795 =>	"00000000",	-- ........
		1796 =>	"00000000",	-- ........
		1797 =>	"00000000",	-- ........
		1798 =>	"11011100",	-- ##.###..
		1799 =>	"01100110",	-- .##..##.
		1800 =>	"01100110",	-- .##..##.
		1801 =>	"01100110",	-- .##..##.
		1802 =>	"01111100",	-- .#####..
		1803 =>	"01100000",	-- .##.....
		1804 =>	"01100000",	-- .##.....
		1805 =>	"11110000",	-- ####....
		1806 =>	"00000000",	-- ........
		1807 =>	"00000000",	-- ........

		-- char 0x71='q'  
		1808 =>	"00000000",	-- ........
		1809 =>	"00000000",	-- ........
		1810 =>	"00000000",	-- ........
		1811 =>	"00000000",	-- ........
		1812 =>	"00000000",	-- ........
		1813 =>	"00000000",	-- ........
		1814 =>	"01110110",	-- .###.##.
		1815 =>	"11001100",	-- ##..##..
		1816 =>	"11001100",	-- ##..##..
		1817 =>	"11001100",	-- ##..##..
		1818 =>	"01111100",	-- .#####..
		1819 =>	"00001100",	-- ....##..
		1820 =>	"00001100",	-- ....##..
		1821 =>	"00011110",	-- ...####.
		1822 =>	"00000000",	-- ........
		1823 =>	"00000000",	-- ........

		-- char 0x72='r'  
		1824 =>	"00000000",	-- ........
		1825 =>	"00000000",	-- ........
		1826 =>	"00000000",	-- ........
		1827 =>	"00000000",	-- ........
		1828 =>	"00000000",	-- ........
		1829 =>	"00000000",	-- ........
		1830 =>	"11011100",	-- ##.###..
		1831 =>	"01110110",	-- .###.##.
		1832 =>	"01100110",	-- .##..##.
		1833 =>	"01100000",	-- .##.....
		1834 =>	"01100000",	-- .##.....
		1835 =>	"11110000",	-- ####....
		1836 =>	"00000000",	-- ........
		1837 =>	"00000000",	-- ........
		1838 =>	"00000000",	-- ........
		1839 =>	"00000000",	-- ........

		-- char 0x73='s'  
		1840 =>	"00000000",	-- ........
		1841 =>	"00000000",	-- ........
		1842 =>	"00000000",	-- ........
		1843 =>	"00000000",	-- ........
		1844 =>	"00000000",	-- ........
		1845 =>	"00000000",	-- ........
		1846 =>	"01111100",	-- .#####..
		1847 =>	"11000110",	-- ##...##.
		1848 =>	"01110000",	-- .###....
		1849 =>	"00011100",	-- ...###..
		1850 =>	"11000110",	-- ##...##.
		1851 =>	"01111100",	-- .#####..
		1852 =>	"00000000",	-- ........
		1853 =>	"00000000",	-- ........
		1854 =>	"00000000",	-- ........
		1855 =>	"00000000",	-- ........

		-- char 0x74='t'  
		1856 =>	"00000000",	-- ........
		1857 =>	"00000000",	-- ........
		1858 =>	"00000000",	-- ........
		1859 =>	"00010000",	-- ...#....
		1860 =>	"00110000",	-- ..##....
		1861 =>	"00110000",	-- ..##....
		1862 =>	"11111100",	-- ######..
		1863 =>	"00110000",	-- ..##....
		1864 =>	"00110000",	-- ..##....
		1865 =>	"00110000",	-- ..##....
		1866 =>	"00110110",	-- ..##.##.
		1867 =>	"00011100",	-- ...###..
		1868 =>	"00000000",	-- ........
		1869 =>	"00000000",	-- ........
		1870 =>	"00000000",	-- ........
		1871 =>	"00000000",	-- ........

		-- char 0x75='u'  
		1872 =>	"00000000",	-- ........
		1873 =>	"00000000",	-- ........
		1874 =>	"00000000",	-- ........
		1875 =>	"00000000",	-- ........
		1876 =>	"00000000",	-- ........
		1877 =>	"00000000",	-- ........
		1878 =>	"11001100",	-- ##..##..
		1879 =>	"11001100",	-- ##..##..
		1880 =>	"11001100",	-- ##..##..
		1881 =>	"11001100",	-- ##..##..
		1882 =>	"11001100",	-- ##..##..
		1883 =>	"01110110",	-- .###.##.
		1884 =>	"00000000",	-- ........
		1885 =>	"00000000",	-- ........
		1886 =>	"00000000",	-- ........
		1887 =>	"00000000",	-- ........

		-- char 0x76='v'  
		1888 =>	"00000000",	-- ........
		1889 =>	"00000000",	-- ........
		1890 =>	"00000000",	-- ........
		1891 =>	"00000000",	-- ........
		1892 =>	"00000000",	-- ........
		1893 =>	"00000000",	-- ........
		1894 =>	"01100110",	-- .##..##.
		1895 =>	"01100110",	-- .##..##.
		1896 =>	"01100110",	-- .##..##.
		1897 =>	"01100110",	-- .##..##.
		1898 =>	"00111100",	-- ..####..
		1899 =>	"00011000",	-- ...##...
		1900 =>	"00000000",	-- ........
		1901 =>	"00000000",	-- ........
		1902 =>	"00000000",	-- ........
		1903 =>	"00000000",	-- ........

		-- char 0x77='w'  
		1904 =>	"00000000",	-- ........
		1905 =>	"00000000",	-- ........
		1906 =>	"00000000",	-- ........
		1907 =>	"00000000",	-- ........
		1908 =>	"00000000",	-- ........
		1909 =>	"00000000",	-- ........
		1910 =>	"11000110",	-- ##...##.
		1911 =>	"11000110",	-- ##...##.
		1912 =>	"11010110",	-- ##.#.##.
		1913 =>	"11010110",	-- ##.#.##.
		1914 =>	"11111110",	-- #######.
		1915 =>	"01101100",	-- .##.##..
		1916 =>	"00000000",	-- ........
		1917 =>	"00000000",	-- ........
		1918 =>	"00000000",	-- ........
		1919 =>	"00000000",	-- ........

		-- char 0x78='x'  
		1920 =>	"00000000",	-- ........
		1921 =>	"00000000",	-- ........
		1922 =>	"00000000",	-- ........
		1923 =>	"00000000",	-- ........
		1924 =>	"00000000",	-- ........
		1925 =>	"00000000",	-- ........
		1926 =>	"11000110",	-- ##...##.
		1927 =>	"01101100",	-- .##.##..
		1928 =>	"00111000",	-- ..###...
		1929 =>	"00111000",	-- ..###...
		1930 =>	"01101100",	-- .##.##..
		1931 =>	"11000110",	-- ##...##.
		1932 =>	"00000000",	-- ........
		1933 =>	"00000000",	-- ........
		1934 =>	"00000000",	-- ........
		1935 =>	"00000000",	-- ........

		-- char 0x79='y'  
		1936 =>	"00000000",	-- ........
		1937 =>	"00000000",	-- ........
		1938 =>	"00000000",	-- ........
		1939 =>	"00000000",	-- ........
		1940 =>	"00000000",	-- ........
		1941 =>	"00000000",	-- ........
		1942 =>	"11000110",	-- ##...##.
		1943 =>	"11000110",	-- ##...##.
		1944 =>	"11000110",	-- ##...##.
		1945 =>	"11000110",	-- ##...##.
		1946 =>	"01111110",	-- .######.
		1947 =>	"00000110",	-- .....##.
		1948 =>	"00001100",	-- ....##..
		1949 =>	"11111000",	-- #####...
		1950 =>	"00000000",	-- ........
		1951 =>	"00000000",	-- ........

		-- char 0x7a='z'  
		1952 =>	"00000000",	-- ........
		1953 =>	"00000000",	-- ........
		1954 =>	"00000000",	-- ........
		1955 =>	"00000000",	-- ........
		1956 =>	"00000000",	-- ........
		1957 =>	"00000000",	-- ........
		1958 =>	"11111110",	-- #######.
		1959 =>	"11001100",	-- ##..##..
		1960 =>	"00011000",	-- ...##...
		1961 =>	"00110000",	-- ..##....
		1962 =>	"01100110",	-- .##..##.
		1963 =>	"11111110",	-- #######.
		1964 =>	"00000000",	-- ........
		1965 =>	"00000000",	-- ........
		1966 =>	"00000000",	-- ........
		1967 =>	"00000000",	-- ........

		-- char 0x7b='{'  
		1968 =>	"00000000",	-- ........
		1969 =>	"00000000",	-- ........
		1970 =>	"00000000",	-- ........
		1971 =>	"00001110",	-- ....###.
		1972 =>	"00011000",	-- ...##...
		1973 =>	"00011000",	-- ...##...
		1974 =>	"00011000",	-- ...##...
		1975 =>	"01110000",	-- .###....
		1976 =>	"00011000",	-- ...##...
		1977 =>	"00011000",	-- ...##...
		1978 =>	"00011000",	-- ...##...
		1979 =>	"00001110",	-- ....###.
		1980 =>	"00000000",	-- ........
		1981 =>	"00000000",	-- ........
		1982 =>	"00000000",	-- ........
		1983 =>	"00000000",	-- ........

		-- char 0x7c='|'  
		1984 =>	"00000000",	-- ........
		1985 =>	"00000000",	-- ........
		1986 =>	"00000000",	-- ........
		1987 =>	"00011000",	-- ...##...
		1988 =>	"00011000",	-- ...##...
		1989 =>	"00011000",	-- ...##...
		1990 =>	"00011000",	-- ...##...
		1991 =>	"00000000",	-- ........
		1992 =>	"00011000",	-- ...##...
		1993 =>	"00011000",	-- ...##...
		1994 =>	"00011000",	-- ...##...
		1995 =>	"00011000",	-- ...##...
		1996 =>	"00000000",	-- ........
		1997 =>	"00000000",	-- ........
		1998 =>	"00000000",	-- ........
		1999 =>	"00000000",	-- ........

		-- char 0x7d='}'  
		2000 =>	"00000000",	-- ........
		2001 =>	"00000000",	-- ........
		2002 =>	"00000000",	-- ........
		2003 =>	"01110000",	-- .###....
		2004 =>	"00011000",	-- ...##...
		2005 =>	"00011000",	-- ...##...
		2006 =>	"00011000",	-- ...##...
		2007 =>	"00001110",	-- ....###.
		2008 =>	"00011000",	-- ...##...
		2009 =>	"00011000",	-- ...##...
		2010 =>	"00011000",	-- ...##...
		2011 =>	"01110000",	-- .###....
		2012 =>	"00000000",	-- ........
		2013 =>	"00000000",	-- ........
		2014 =>	"00000000",	-- ........
		2015 =>	"00000000",	-- ........

		-- char 0x7e='~'  
		2016 =>	"00000000",	-- ........
		2017 =>	"00000000",	-- ........
		2018 =>	"00000000",	-- ........
		2019 =>	"01110110",	-- .###.##.
		2020 =>	"11011100",	-- ##.###..
		2021 =>	"00000000",	-- ........
		2022 =>	"00000000",	-- ........
		2023 =>	"00000000",	-- ........
		2024 =>	"00000000",	-- ........
		2025 =>	"00000000",	-- ........
		2026 =>	"00000000",	-- ........
		2027 =>	"00000000",	-- ........
		2028 =>	"00000000",	-- ........
		2029 =>	"00000000",	-- ........
		2030 =>	"00000000",	-- ........
		2031 =>	"00000000",	-- ........

		-- char 0x7f='\x7f
		2032 =>	"00000000",	-- ........
		2033 =>	"00000000",	-- ........
		2034 =>	"00000000",	-- ........
		2035 =>	"00000000",	-- ........
		2036 =>	"00000000",	-- ........
		2037 =>	"00010000",	-- ...#....
		2038 =>	"00111000",	-- ..###...
		2039 =>	"01101100",	-- .##.##..
		2040 =>	"11000110",	-- ##...##.
		2041 =>	"11000110",	-- ##...##.
		2042 =>	"11111110",	-- #######.
		2043 =>	"00000000",	-- ........
		2044 =>	"00000000",	-- ........
		2045 =>	"00000000",	-- ........
		2046 =>	"00000000",	-- ........
		2047 =>	"00000000",	-- ........

		-- char 0x80='\x80
		2048 =>	"00000000",	-- ........
		2049 =>	"00000000",	-- ........
		2050 =>	"00000000",	-- ........
		2051 =>	"00111100",	-- ..####..
		2052 =>	"01100110",	-- .##..##.
		2053 =>	"11000010",	-- ##....#.
		2054 =>	"11000000",	-- ##......
		2055 =>	"11000000",	-- ##......
		2056 =>	"11000010",	-- ##....#.
		2057 =>	"01100110",	-- .##..##.
		2058 =>	"00111100",	-- ..####..
		2059 =>	"00001100",	-- ....##..
		2060 =>	"00000110",	-- .....##.
		2061 =>	"01111100",	-- .#####..
		2062 =>	"00000000",	-- ........
		2063 =>	"00000000",	-- ........

		-- char 0x81='\x81
		2064 =>	"00000000",	-- ........
		2065 =>	"00000000",	-- ........
		2066 =>	"00000000",	-- ........
		2067 =>	"11001100",	-- ##..##..
		2068 =>	"11001100",	-- ##..##..
		2069 =>	"00000000",	-- ........
		2070 =>	"11001100",	-- ##..##..
		2071 =>	"11001100",	-- ##..##..
		2072 =>	"11001100",	-- ##..##..
		2073 =>	"11001100",	-- ##..##..
		2074 =>	"11001100",	-- ##..##..
		2075 =>	"01110110",	-- .###.##.
		2076 =>	"00000000",	-- ........
		2077 =>	"00000000",	-- ........
		2078 =>	"00000000",	-- ........
		2079 =>	"00000000",	-- ........

		-- char 0x82='\x82
		2080 =>	"00000000",	-- ........
		2081 =>	"00000000",	-- ........
		2082 =>	"00001100",	-- ....##..
		2083 =>	"00011000",	-- ...##...
		2084 =>	"00110000",	-- ..##....
		2085 =>	"00000000",	-- ........
		2086 =>	"01111100",	-- .#####..
		2087 =>	"11000110",	-- ##...##.
		2088 =>	"11111110",	-- #######.
		2089 =>	"11000000",	-- ##......
		2090 =>	"11000110",	-- ##...##.
		2091 =>	"01111100",	-- .#####..
		2092 =>	"00000000",	-- ........
		2093 =>	"00000000",	-- ........
		2094 =>	"00000000",	-- ........
		2095 =>	"00000000",	-- ........

		-- char 0x83='\x83
		2096 =>	"00000000",	-- ........
		2097 =>	"00000000",	-- ........
		2098 =>	"00010000",	-- ...#....
		2099 =>	"00111000",	-- ..###...
		2100 =>	"01101100",	-- .##.##..
		2101 =>	"00000000",	-- ........
		2102 =>	"01111000",	-- .####...
		2103 =>	"00001100",	-- ....##..
		2104 =>	"01111100",	-- .#####..
		2105 =>	"11001100",	-- ##..##..
		2106 =>	"11001100",	-- ##..##..
		2107 =>	"01110110",	-- .###.##.
		2108 =>	"00000000",	-- ........
		2109 =>	"00000000",	-- ........
		2110 =>	"00000000",	-- ........
		2111 =>	"00000000",	-- ........

		-- char 0x84='\x84
		2112 =>	"00000000",	-- ........
		2113 =>	"00000000",	-- ........
		2114 =>	"00000000",	-- ........
		2115 =>	"11001100",	-- ##..##..
		2116 =>	"11001100",	-- ##..##..
		2117 =>	"00000000",	-- ........
		2118 =>	"01111000",	-- .####...
		2119 =>	"00001100",	-- ....##..
		2120 =>	"01111100",	-- .#####..
		2121 =>	"11001100",	-- ##..##..
		2122 =>	"11001100",	-- ##..##..
		2123 =>	"01110110",	-- .###.##.
		2124 =>	"00000000",	-- ........
		2125 =>	"00000000",	-- ........
		2126 =>	"00000000",	-- ........
		2127 =>	"00000000",	-- ........

		-- char 0x85='\x85
		2128 =>	"00000000",	-- ........
		2129 =>	"00000000",	-- ........
		2130 =>	"01100000",	-- .##.....
		2131 =>	"00110000",	-- ..##....
		2132 =>	"00011000",	-- ...##...
		2133 =>	"00000000",	-- ........
		2134 =>	"01111000",	-- .####...
		2135 =>	"00001100",	-- ....##..
		2136 =>	"01111100",	-- .#####..
		2137 =>	"11001100",	-- ##..##..
		2138 =>	"11001100",	-- ##..##..
		2139 =>	"01110110",	-- .###.##.
		2140 =>	"00000000",	-- ........
		2141 =>	"00000000",	-- ........
		2142 =>	"00000000",	-- ........
		2143 =>	"00000000",	-- ........

		-- char 0x86='\x86
		2144 =>	"00000000",	-- ........
		2145 =>	"00000000",	-- ........
		2146 =>	"00111000",	-- ..###...
		2147 =>	"01101100",	-- .##.##..
		2148 =>	"00111000",	-- ..###...
		2149 =>	"00000000",	-- ........
		2150 =>	"01111000",	-- .####...
		2151 =>	"00001100",	-- ....##..
		2152 =>	"01111100",	-- .#####..
		2153 =>	"11001100",	-- ##..##..
		2154 =>	"11001100",	-- ##..##..
		2155 =>	"01110110",	-- .###.##.
		2156 =>	"00000000",	-- ........
		2157 =>	"00000000",	-- ........
		2158 =>	"00000000",	-- ........
		2159 =>	"00000000",	-- ........

		-- char 0x87='\x87
		2160 =>	"00000000",	-- ........
		2161 =>	"00000000",	-- ........
		2162 =>	"00000000",	-- ........
		2163 =>	"00000000",	-- ........
		2164 =>	"00000000",	-- ........
		2165 =>	"00111100",	-- ..####..
		2166 =>	"01100110",	-- .##..##.
		2167 =>	"01100000",	-- .##.....
		2168 =>	"01100110",	-- .##..##.
		2169 =>	"00111100",	-- ..####..
		2170 =>	"00001100",	-- ....##..
		2171 =>	"00000110",	-- .....##.
		2172 =>	"00111100",	-- ..####..
		2173 =>	"00000000",	-- ........
		2174 =>	"00000000",	-- ........
		2175 =>	"00000000",	-- ........

		-- char 0x88='\x88
		2176 =>	"00000000",	-- ........
		2177 =>	"00000000",	-- ........
		2178 =>	"00010000",	-- ...#....
		2179 =>	"00111000",	-- ..###...
		2180 =>	"01101100",	-- .##.##..
		2181 =>	"00000000",	-- ........
		2182 =>	"01111100",	-- .#####..
		2183 =>	"11000110",	-- ##...##.
		2184 =>	"11111110",	-- #######.
		2185 =>	"11000000",	-- ##......
		2186 =>	"11000110",	-- ##...##.
		2187 =>	"01111100",	-- .#####..
		2188 =>	"00000000",	-- ........
		2189 =>	"00000000",	-- ........
		2190 =>	"00000000",	-- ........
		2191 =>	"00000000",	-- ........

		-- char 0x89='\x89
		2192 =>	"00000000",	-- ........
		2193 =>	"00000000",	-- ........
		2194 =>	"00000000",	-- ........
		2195 =>	"11001100",	-- ##..##..
		2196 =>	"11001100",	-- ##..##..
		2197 =>	"00000000",	-- ........
		2198 =>	"01111100",	-- .#####..
		2199 =>	"11000110",	-- ##...##.
		2200 =>	"11111110",	-- #######.
		2201 =>	"11000000",	-- ##......
		2202 =>	"11000110",	-- ##...##.
		2203 =>	"01111100",	-- .#####..
		2204 =>	"00000000",	-- ........
		2205 =>	"00000000",	-- ........
		2206 =>	"00000000",	-- ........
		2207 =>	"00000000",	-- ........

		-- char 0x8a='\x8a
		2208 =>	"00000000",	-- ........
		2209 =>	"00000000",	-- ........
		2210 =>	"01100000",	-- .##.....
		2211 =>	"00110000",	-- ..##....
		2212 =>	"00011000",	-- ...##...
		2213 =>	"00000000",	-- ........
		2214 =>	"01111100",	-- .#####..
		2215 =>	"11000110",	-- ##...##.
		2216 =>	"11111110",	-- #######.
		2217 =>	"11000000",	-- ##......
		2218 =>	"11000110",	-- ##...##.
		2219 =>	"01111100",	-- .#####..
		2220 =>	"00000000",	-- ........
		2221 =>	"00000000",	-- ........
		2222 =>	"00000000",	-- ........
		2223 =>	"00000000",	-- ........

		-- char 0x8b='\x8b
		2224 =>	"00000000",	-- ........
		2225 =>	"00000000",	-- ........
		2226 =>	"00000000",	-- ........
		2227 =>	"01100110",	-- .##..##.
		2228 =>	"01100110",	-- .##..##.
		2229 =>	"00000000",	-- ........
		2230 =>	"00111000",	-- ..###...
		2231 =>	"00011000",	-- ...##...
		2232 =>	"00011000",	-- ...##...
		2233 =>	"00011000",	-- ...##...
		2234 =>	"00011000",	-- ...##...
		2235 =>	"00111100",	-- ..####..
		2236 =>	"00000000",	-- ........
		2237 =>	"00000000",	-- ........
		2238 =>	"00000000",	-- ........
		2239 =>	"00000000",	-- ........

		-- char 0x8c='\x8c
		2240 =>	"00000000",	-- ........
		2241 =>	"00000000",	-- ........
		2242 =>	"00011000",	-- ...##...
		2243 =>	"00111100",	-- ..####..
		2244 =>	"01100110",	-- .##..##.
		2245 =>	"00000000",	-- ........
		2246 =>	"00111000",	-- ..###...
		2247 =>	"00011000",	-- ...##...
		2248 =>	"00011000",	-- ...##...
		2249 =>	"00011000",	-- ...##...
		2250 =>	"00011000",	-- ...##...
		2251 =>	"00111100",	-- ..####..
		2252 =>	"00000000",	-- ........
		2253 =>	"00000000",	-- ........
		2254 =>	"00000000",	-- ........
		2255 =>	"00000000",	-- ........

		-- char 0x8d='\x8d
		2256 =>	"00000000",	-- ........
		2257 =>	"00000000",	-- ........
		2258 =>	"01100000",	-- .##.....
		2259 =>	"00110000",	-- ..##....
		2260 =>	"00011000",	-- ...##...
		2261 =>	"00000000",	-- ........
		2262 =>	"00111000",	-- ..###...
		2263 =>	"00011000",	-- ...##...
		2264 =>	"00011000",	-- ...##...
		2265 =>	"00011000",	-- ...##...
		2266 =>	"00011000",	-- ...##...
		2267 =>	"00111100",	-- ..####..
		2268 =>	"00000000",	-- ........
		2269 =>	"00000000",	-- ........
		2270 =>	"00000000",	-- ........
		2271 =>	"00000000",	-- ........

		-- char 0x8e='\x8e
		2272 =>	"00000000",	-- ........
		2273 =>	"00000000",	-- ........
		2274 =>	"11000110",	-- ##...##.
		2275 =>	"11000110",	-- ##...##.
		2276 =>	"00010000",	-- ...#....
		2277 =>	"00111000",	-- ..###...
		2278 =>	"01101100",	-- .##.##..
		2279 =>	"11000110",	-- ##...##.
		2280 =>	"11000110",	-- ##...##.
		2281 =>	"11111110",	-- #######.
		2282 =>	"11000110",	-- ##...##.
		2283 =>	"11000110",	-- ##...##.
		2284 =>	"00000000",	-- ........
		2285 =>	"00000000",	-- ........
		2286 =>	"00000000",	-- ........
		2287 =>	"00000000",	-- ........

		-- char 0x8f='\x8f
		2288 =>	"00000000",	-- ........
		2289 =>	"00111000",	-- ..###...
		2290 =>	"01101100",	-- .##.##..
		2291 =>	"00111000",	-- ..###...
		2292 =>	"00000000",	-- ........
		2293 =>	"00111000",	-- ..###...
		2294 =>	"01101100",	-- .##.##..
		2295 =>	"11000110",	-- ##...##.
		2296 =>	"11000110",	-- ##...##.
		2297 =>	"11111110",	-- #######.
		2298 =>	"11000110",	-- ##...##.
		2299 =>	"11000110",	-- ##...##.
		2300 =>	"00000000",	-- ........
		2301 =>	"00000000",	-- ........
		2302 =>	"00000000",	-- ........
		2303 =>	"00000000",	-- ........

		-- char 0x90='\x90
		2304 =>	"00000000",	-- ........
		2305 =>	"00011000",	-- ...##...
		2306 =>	"00110000",	-- ..##....
		2307 =>	"01100000",	-- .##.....
		2308 =>	"00000000",	-- ........
		2309 =>	"11111110",	-- #######.
		2310 =>	"01100110",	-- .##..##.
		2311 =>	"01100000",	-- .##.....
		2312 =>	"01111100",	-- .#####..
		2313 =>	"01100000",	-- .##.....
		2314 =>	"01100110",	-- .##..##.
		2315 =>	"11111110",	-- #######.
		2316 =>	"00000000",	-- ........
		2317 =>	"00000000",	-- ........
		2318 =>	"00000000",	-- ........
		2319 =>	"00000000",	-- ........

		-- char 0x91='\x91
		2320 =>	"00000000",	-- ........
		2321 =>	"00000000",	-- ........
		2322 =>	"00000000",	-- ........
		2323 =>	"00000000",	-- ........
		2324 =>	"00000000",	-- ........
		2325 =>	"11001100",	-- ##..##..
		2326 =>	"01110110",	-- .###.##.
		2327 =>	"00110110",	-- ..##.##.
		2328 =>	"01111110",	-- .######.
		2329 =>	"11011000",	-- ##.##...
		2330 =>	"11011000",	-- ##.##...
		2331 =>	"01101110",	-- .##.###.
		2332 =>	"00000000",	-- ........
		2333 =>	"00000000",	-- ........
		2334 =>	"00000000",	-- ........
		2335 =>	"00000000",	-- ........

		-- char 0x92='\x92
		2336 =>	"00000000",	-- ........
		2337 =>	"00000000",	-- ........
		2338 =>	"00000000",	-- ........
		2339 =>	"00111110",	-- ..#####.
		2340 =>	"01101100",	-- .##.##..
		2341 =>	"11001100",	-- ##..##..
		2342 =>	"11001100",	-- ##..##..
		2343 =>	"11111110",	-- #######.
		2344 =>	"11001100",	-- ##..##..
		2345 =>	"11001100",	-- ##..##..
		2346 =>	"11001100",	-- ##..##..
		2347 =>	"11001110",	-- ##..###.
		2348 =>	"00000000",	-- ........
		2349 =>	"00000000",	-- ........
		2350 =>	"00000000",	-- ........
		2351 =>	"00000000",	-- ........

		-- char 0x93='\x93
		2352 =>	"00000000",	-- ........
		2353 =>	"00000000",	-- ........
		2354 =>	"00010000",	-- ...#....
		2355 =>	"00111000",	-- ..###...
		2356 =>	"01101100",	-- .##.##..
		2357 =>	"00000000",	-- ........
		2358 =>	"01111100",	-- .#####..
		2359 =>	"11000110",	-- ##...##.
		2360 =>	"11000110",	-- ##...##.
		2361 =>	"11000110",	-- ##...##.
		2362 =>	"11000110",	-- ##...##.
		2363 =>	"01111100",	-- .#####..
		2364 =>	"00000000",	-- ........
		2365 =>	"00000000",	-- ........
		2366 =>	"00000000",	-- ........
		2367 =>	"00000000",	-- ........

		-- char 0x94='\x94
		2368 =>	"00000000",	-- ........
		2369 =>	"00000000",	-- ........
		2370 =>	"00000000",	-- ........
		2371 =>	"11000110",	-- ##...##.
		2372 =>	"11000110",	-- ##...##.
		2373 =>	"00000000",	-- ........
		2374 =>	"01111100",	-- .#####..
		2375 =>	"11000110",	-- ##...##.
		2376 =>	"11000110",	-- ##...##.
		2377 =>	"11000110",	-- ##...##.
		2378 =>	"11000110",	-- ##...##.
		2379 =>	"01111100",	-- .#####..
		2380 =>	"00000000",	-- ........
		2381 =>	"00000000",	-- ........
		2382 =>	"00000000",	-- ........
		2383 =>	"00000000",	-- ........

		-- char 0x95='\x95
		2384 =>	"00000000",	-- ........
		2385 =>	"00000000",	-- ........
		2386 =>	"01100000",	-- .##.....
		2387 =>	"00110000",	-- ..##....
		2388 =>	"00011000",	-- ...##...
		2389 =>	"00000000",	-- ........
		2390 =>	"01111100",	-- .#####..
		2391 =>	"11000110",	-- ##...##.
		2392 =>	"11000110",	-- ##...##.
		2393 =>	"11000110",	-- ##...##.
		2394 =>	"11000110",	-- ##...##.
		2395 =>	"01111100",	-- .#####..
		2396 =>	"00000000",	-- ........
		2397 =>	"00000000",	-- ........
		2398 =>	"00000000",	-- ........
		2399 =>	"00000000",	-- ........

		-- char 0x96='\x96
		2400 =>	"00000000",	-- ........
		2401 =>	"00000000",	-- ........
		2402 =>	"00110000",	-- ..##....
		2403 =>	"01111000",	-- .####...
		2404 =>	"11001100",	-- ##..##..
		2405 =>	"00000000",	-- ........
		2406 =>	"11001100",	-- ##..##..
		2407 =>	"11001100",	-- ##..##..
		2408 =>	"11001100",	-- ##..##..
		2409 =>	"11001100",	-- ##..##..
		2410 =>	"11001100",	-- ##..##..
		2411 =>	"01110110",	-- .###.##.
		2412 =>	"00000000",	-- ........
		2413 =>	"00000000",	-- ........
		2414 =>	"00000000",	-- ........
		2415 =>	"00000000",	-- ........

		-- char 0x97='\x97
		2416 =>	"00000000",	-- ........
		2417 =>	"00000000",	-- ........
		2418 =>	"01100000",	-- .##.....
		2419 =>	"00110000",	-- ..##....
		2420 =>	"00011000",	-- ...##...
		2421 =>	"00000000",	-- ........
		2422 =>	"11001100",	-- ##..##..
		2423 =>	"11001100",	-- ##..##..
		2424 =>	"11001100",	-- ##..##..
		2425 =>	"11001100",	-- ##..##..
		2426 =>	"11001100",	-- ##..##..
		2427 =>	"01110110",	-- .###.##.
		2428 =>	"00000000",	-- ........
		2429 =>	"00000000",	-- ........
		2430 =>	"00000000",	-- ........
		2431 =>	"00000000",	-- ........

		-- char 0x98='\x98
		2432 =>	"00000000",	-- ........
		2433 =>	"00000000",	-- ........
		2434 =>	"00000000",	-- ........
		2435 =>	"11000110",	-- ##...##.
		2436 =>	"11000110",	-- ##...##.
		2437 =>	"00000000",	-- ........
		2438 =>	"11000110",	-- ##...##.
		2439 =>	"11000110",	-- ##...##.
		2440 =>	"11000110",	-- ##...##.
		2441 =>	"11000110",	-- ##...##.
		2442 =>	"01111110",	-- .######.
		2443 =>	"00000110",	-- .....##.
		2444 =>	"00001100",	-- ....##..
		2445 =>	"01111000",	-- .####...
		2446 =>	"00000000",	-- ........
		2447 =>	"00000000",	-- ........

		-- char 0x99='\x99
		2448 =>	"00000000",	-- ........
		2449 =>	"00000000",	-- ........
		2450 =>	"11000110",	-- ##...##.
		2451 =>	"11000110",	-- ##...##.
		2452 =>	"00111000",	-- ..###...
		2453 =>	"01101100",	-- .##.##..
		2454 =>	"11000110",	-- ##...##.
		2455 =>	"11000110",	-- ##...##.
		2456 =>	"11000110",	-- ##...##.
		2457 =>	"11000110",	-- ##...##.
		2458 =>	"01101100",	-- .##.##..
		2459 =>	"00111000",	-- ..###...
		2460 =>	"00000000",	-- ........
		2461 =>	"00000000",	-- ........
		2462 =>	"00000000",	-- ........
		2463 =>	"00000000",	-- ........

		-- char 0x9a='\x9a
		2464 =>	"00000000",	-- ........
		2465 =>	"00000000",	-- ........
		2466 =>	"11000110",	-- ##...##.
		2467 =>	"11000110",	-- ##...##.
		2468 =>	"00000000",	-- ........
		2469 =>	"11000110",	-- ##...##.
		2470 =>	"11000110",	-- ##...##.
		2471 =>	"11000110",	-- ##...##.
		2472 =>	"11000110",	-- ##...##.
		2473 =>	"11000110",	-- ##...##.
		2474 =>	"11000110",	-- ##...##.
		2475 =>	"01111100",	-- .#####..
		2476 =>	"00000000",	-- ........
		2477 =>	"00000000",	-- ........
		2478 =>	"00000000",	-- ........
		2479 =>	"00000000",	-- ........

		-- char 0x9b='\x9b
		2480 =>	"00000000",	-- ........
		2481 =>	"00000000",	-- ........
		2482 =>	"00011000",	-- ...##...
		2483 =>	"00011000",	-- ...##...
		2484 =>	"00111100",	-- ..####..
		2485 =>	"01100110",	-- .##..##.
		2486 =>	"01100000",	-- .##.....
		2487 =>	"01100000",	-- .##.....
		2488 =>	"01100110",	-- .##..##.
		2489 =>	"00111100",	-- ..####..
		2490 =>	"00011000",	-- ...##...
		2491 =>	"00011000",	-- ...##...
		2492 =>	"00000000",	-- ........
		2493 =>	"00000000",	-- ........
		2494 =>	"00000000",	-- ........
		2495 =>	"00000000",	-- ........

		-- char 0x9c='\x9c
		2496 =>	"00000000",	-- ........
		2497 =>	"00000000",	-- ........
		2498 =>	"00111000",	-- ..###...
		2499 =>	"01101100",	-- .##.##..
		2500 =>	"01100100",	-- .##..#..
		2501 =>	"01100000",	-- .##.....
		2502 =>	"11110000",	-- ####....
		2503 =>	"01100000",	-- .##.....
		2504 =>	"01100000",	-- .##.....
		2505 =>	"01100000",	-- .##.....
		2506 =>	"11100110",	-- ###..##.
		2507 =>	"11111100",	-- ######..
		2508 =>	"00000000",	-- ........
		2509 =>	"00000000",	-- ........
		2510 =>	"00000000",	-- ........
		2511 =>	"00000000",	-- ........

		-- char 0x9d='\x9d
		2512 =>	"00000000",	-- ........
		2513 =>	"00000000",	-- ........
		2514 =>	"00000000",	-- ........
		2515 =>	"01100110",	-- .##..##.
		2516 =>	"01100110",	-- .##..##.
		2517 =>	"00111100",	-- ..####..
		2518 =>	"00011000",	-- ...##...
		2519 =>	"01111110",	-- .######.
		2520 =>	"00011000",	-- ...##...
		2521 =>	"01111110",	-- .######.
		2522 =>	"00011000",	-- ...##...
		2523 =>	"00011000",	-- ...##...
		2524 =>	"00000000",	-- ........
		2525 =>	"00000000",	-- ........
		2526 =>	"00000000",	-- ........
		2527 =>	"00000000",	-- ........

		-- char 0x9e='\x9e
		2528 =>	"00000000",	-- ........
		2529 =>	"00000000",	-- ........
		2530 =>	"11111000",	-- #####...
		2531 =>	"11001100",	-- ##..##..
		2532 =>	"11001100",	-- ##..##..
		2533 =>	"11111000",	-- #####...
		2534 =>	"11000100",	-- ##...#..
		2535 =>	"11001100",	-- ##..##..
		2536 =>	"11011110",	-- ##.####.
		2537 =>	"11001100",	-- ##..##..
		2538 =>	"11001100",	-- ##..##..
		2539 =>	"11000110",	-- ##...##.
		2540 =>	"00000000",	-- ........
		2541 =>	"00000000",	-- ........
		2542 =>	"00000000",	-- ........
		2543 =>	"00000000",	-- ........

		-- char 0x9f='\x9f
		2544 =>	"00000000",	-- ........
		2545 =>	"00000000",	-- ........
		2546 =>	"00001110",	-- ....###.
		2547 =>	"00011011",	-- ...##.##
		2548 =>	"00011000",	-- ...##...
		2549 =>	"00011000",	-- ...##...
		2550 =>	"00011000",	-- ...##...
		2551 =>	"01111110",	-- .######.
		2552 =>	"00011000",	-- ...##...
		2553 =>	"00011000",	-- ...##...
		2554 =>	"00011000",	-- ...##...
		2555 =>	"00011000",	-- ...##...
		2556 =>	"11011000",	-- ##.##...
		2557 =>	"01110000",	-- .###....
		2558 =>	"00000000",	-- ........
		2559 =>	"00000000",	-- ........

		-- char 0xa0='\xa0
		2560 =>	"00000000",	-- ........
		2561 =>	"00000000",	-- ........
		2562 =>	"00011000",	-- ...##...
		2563 =>	"00110000",	-- ..##....
		2564 =>	"01100000",	-- .##.....
		2565 =>	"00000000",	-- ........
		2566 =>	"01111000",	-- .####...
		2567 =>	"00001100",	-- ....##..
		2568 =>	"01111100",	-- .#####..
		2569 =>	"11001100",	-- ##..##..
		2570 =>	"11001100",	-- ##..##..
		2571 =>	"01110110",	-- .###.##.
		2572 =>	"00000000",	-- ........
		2573 =>	"00000000",	-- ........
		2574 =>	"00000000",	-- ........
		2575 =>	"00000000",	-- ........

		-- char 0xa1='\xa1
		2576 =>	"00000000",	-- ........
		2577 =>	"00000000",	-- ........
		2578 =>	"00001100",	-- ....##..
		2579 =>	"00011000",	-- ...##...
		2580 =>	"00110000",	-- ..##....
		2581 =>	"00000000",	-- ........
		2582 =>	"00111000",	-- ..###...
		2583 =>	"00011000",	-- ...##...
		2584 =>	"00011000",	-- ...##...
		2585 =>	"00011000",	-- ...##...
		2586 =>	"00011000",	-- ...##...
		2587 =>	"00111100",	-- ..####..
		2588 =>	"00000000",	-- ........
		2589 =>	"00000000",	-- ........
		2590 =>	"00000000",	-- ........
		2591 =>	"00000000",	-- ........

		-- char 0xa2='\xa2
		2592 =>	"00000000",	-- ........
		2593 =>	"00000000",	-- ........
		2594 =>	"00011000",	-- ...##...
		2595 =>	"00110000",	-- ..##....
		2596 =>	"01100000",	-- .##.....
		2597 =>	"00000000",	-- ........
		2598 =>	"01111100",	-- .#####..
		2599 =>	"11000110",	-- ##...##.
		2600 =>	"11000110",	-- ##...##.
		2601 =>	"11000110",	-- ##...##.
		2602 =>	"11000110",	-- ##...##.
		2603 =>	"01111100",	-- .#####..
		2604 =>	"00000000",	-- ........
		2605 =>	"00000000",	-- ........
		2606 =>	"00000000",	-- ........
		2607 =>	"00000000",	-- ........

		-- char 0xa3='\xa3
		2608 =>	"00000000",	-- ........
		2609 =>	"00000000",	-- ........
		2610 =>	"00011000",	-- ...##...
		2611 =>	"00110000",	-- ..##....
		2612 =>	"01100000",	-- .##.....
		2613 =>	"00000000",	-- ........
		2614 =>	"11001100",	-- ##..##..
		2615 =>	"11001100",	-- ##..##..
		2616 =>	"11001100",	-- ##..##..
		2617 =>	"11001100",	-- ##..##..
		2618 =>	"11001100",	-- ##..##..
		2619 =>	"01110110",	-- .###.##.
		2620 =>	"00000000",	-- ........
		2621 =>	"00000000",	-- ........
		2622 =>	"00000000",	-- ........
		2623 =>	"00000000",	-- ........

		-- char 0xa4='\xa4
		2624 =>	"00000000",	-- ........
		2625 =>	"00000000",	-- ........
		2626 =>	"00000000",	-- ........
		2627 =>	"01110110",	-- .###.##.
		2628 =>	"11011100",	-- ##.###..
		2629 =>	"00000000",	-- ........
		2630 =>	"11011100",	-- ##.###..
		2631 =>	"01100110",	-- .##..##.
		2632 =>	"01100110",	-- .##..##.
		2633 =>	"01100110",	-- .##..##.
		2634 =>	"01100110",	-- .##..##.
		2635 =>	"01100110",	-- .##..##.
		2636 =>	"00000000",	-- ........
		2637 =>	"00000000",	-- ........
		2638 =>	"00000000",	-- ........
		2639 =>	"00000000",	-- ........

		-- char 0xa5='\xa5
		2640 =>	"00000000",	-- ........
		2641 =>	"01110110",	-- .###.##.
		2642 =>	"11011100",	-- ##.###..
		2643 =>	"00000000",	-- ........
		2644 =>	"11000110",	-- ##...##.
		2645 =>	"11100110",	-- ###..##.
		2646 =>	"11110110",	-- ####.##.
		2647 =>	"11111110",	-- #######.
		2648 =>	"11011110",	-- ##.####.
		2649 =>	"11001110",	-- ##..###.
		2650 =>	"11000110",	-- ##...##.
		2651 =>	"11000110",	-- ##...##.
		2652 =>	"00000000",	-- ........
		2653 =>	"00000000",	-- ........
		2654 =>	"00000000",	-- ........
		2655 =>	"00000000",	-- ........

		-- char 0xa6='\xa6
		2656 =>	"00000000",	-- ........
		2657 =>	"00000000",	-- ........
		2658 =>	"00111100",	-- ..####..
		2659 =>	"01101100",	-- .##.##..
		2660 =>	"01101100",	-- .##.##..
		2661 =>	"00111110",	-- ..#####.
		2662 =>	"00000000",	-- ........
		2663 =>	"01111110",	-- .######.
		2664 =>	"00000000",	-- ........
		2665 =>	"00000000",	-- ........
		2666 =>	"00000000",	-- ........
		2667 =>	"00000000",	-- ........
		2668 =>	"00000000",	-- ........
		2669 =>	"00000000",	-- ........
		2670 =>	"00000000",	-- ........
		2671 =>	"00000000",	-- ........

		-- char 0xa7='\xa7
		2672 =>	"00000000",	-- ........
		2673 =>	"00000000",	-- ........
		2674 =>	"00111000",	-- ..###...
		2675 =>	"01101100",	-- .##.##..
		2676 =>	"01101100",	-- .##.##..
		2677 =>	"00111000",	-- ..###...
		2678 =>	"00000000",	-- ........
		2679 =>	"01111100",	-- .#####..
		2680 =>	"00000000",	-- ........
		2681 =>	"00000000",	-- ........
		2682 =>	"00000000",	-- ........
		2683 =>	"00000000",	-- ........
		2684 =>	"00000000",	-- ........
		2685 =>	"00000000",	-- ........
		2686 =>	"00000000",	-- ........
		2687 =>	"00000000",	-- ........

		-- char 0xa8='\xa8
		2688 =>	"00000000",	-- ........
		2689 =>	"00000000",	-- ........
		2690 =>	"00000000",	-- ........
		2691 =>	"00110000",	-- ..##....
		2692 =>	"00110000",	-- ..##....
		2693 =>	"00000000",	-- ........
		2694 =>	"00110000",	-- ..##....
		2695 =>	"00110000",	-- ..##....
		2696 =>	"01100000",	-- .##.....
		2697 =>	"11000110",	-- ##...##.
		2698 =>	"11000110",	-- ##...##.
		2699 =>	"01111100",	-- .#####..
		2700 =>	"00000000",	-- ........
		2701 =>	"00000000",	-- ........
		2702 =>	"00000000",	-- ........
		2703 =>	"00000000",	-- ........

		-- char 0xa9='\xa9
		2704 =>	"00000000",	-- ........
		2705 =>	"00000000",	-- ........
		2706 =>	"00000000",	-- ........
		2707 =>	"00000000",	-- ........
		2708 =>	"00000000",	-- ........
		2709 =>	"00000000",	-- ........
		2710 =>	"00000000",	-- ........
		2711 =>	"11111110",	-- #######.
		2712 =>	"11000000",	-- ##......
		2713 =>	"11000000",	-- ##......
		2714 =>	"11000000",	-- ##......
		2715 =>	"00000000",	-- ........
		2716 =>	"00000000",	-- ........
		2717 =>	"00000000",	-- ........
		2718 =>	"00000000",	-- ........
		2719 =>	"00000000",	-- ........

		-- char 0xaa='\xaa
		2720 =>	"00000000",	-- ........
		2721 =>	"00000000",	-- ........
		2722 =>	"00000000",	-- ........
		2723 =>	"00000000",	-- ........
		2724 =>	"00000000",	-- ........
		2725 =>	"00000000",	-- ........
		2726 =>	"00000000",	-- ........
		2727 =>	"11111110",	-- #######.
		2728 =>	"00000110",	-- .....##.
		2729 =>	"00000110",	-- .....##.
		2730 =>	"00000110",	-- .....##.
		2731 =>	"00000000",	-- ........
		2732 =>	"00000000",	-- ........
		2733 =>	"00000000",	-- ........
		2734 =>	"00000000",	-- ........
		2735 =>	"00000000",	-- ........

		-- char 0xab='\xab
		2736 =>	"00000000",	-- ........
		2737 =>	"00000000",	-- ........
		2738 =>	"11000000",	-- ##......
		2739 =>	"11000000",	-- ##......
		2740 =>	"11000110",	-- ##...##.
		2741 =>	"11001100",	-- ##..##..
		2742 =>	"11011000",	-- ##.##...
		2743 =>	"00110000",	-- ..##....
		2744 =>	"01100000",	-- .##.....
		2745 =>	"11011100",	-- ##.###..
		2746 =>	"10000110",	-- #....##.
		2747 =>	"00001100",	-- ....##..
		2748 =>	"00011000",	-- ...##...
		2749 =>	"00111110",	-- ..#####.
		2750 =>	"00000000",	-- ........
		2751 =>	"00000000",	-- ........

		-- char 0xac='\xac
		2752 =>	"00000000",	-- ........
		2753 =>	"00000000",	-- ........
		2754 =>	"11000000",	-- ##......
		2755 =>	"11000000",	-- ##......
		2756 =>	"11000110",	-- ##...##.
		2757 =>	"11001100",	-- ##..##..
		2758 =>	"11011000",	-- ##.##...
		2759 =>	"00110000",	-- ..##....
		2760 =>	"01100110",	-- .##..##.
		2761 =>	"11001110",	-- ##..###.
		2762 =>	"10011110",	-- #..####.
		2763 =>	"00111110",	-- ..#####.
		2764 =>	"00000110",	-- .....##.
		2765 =>	"00000110",	-- .....##.
		2766 =>	"00000000",	-- ........
		2767 =>	"00000000",	-- ........

		-- char 0xad='\xad
		2768 =>	"00000000",	-- ........
		2769 =>	"00000000",	-- ........
		2770 =>	"00000000",	-- ........
		2771 =>	"00011000",	-- ...##...
		2772 =>	"00011000",	-- ...##...
		2773 =>	"00000000",	-- ........
		2774 =>	"00011000",	-- ...##...
		2775 =>	"00011000",	-- ...##...
		2776 =>	"00111100",	-- ..####..
		2777 =>	"00111100",	-- ..####..
		2778 =>	"00111100",	-- ..####..
		2779 =>	"00011000",	-- ...##...
		2780 =>	"00000000",	-- ........
		2781 =>	"00000000",	-- ........
		2782 =>	"00000000",	-- ........
		2783 =>	"00000000",	-- ........

		-- char 0xae='\xae
		2784 =>	"00000000",	-- ........
		2785 =>	"00000000",	-- ........
		2786 =>	"00000000",	-- ........
		2787 =>	"00000000",	-- ........
		2788 =>	"00000000",	-- ........
		2789 =>	"00110110",	-- ..##.##.
		2790 =>	"01101100",	-- .##.##..
		2791 =>	"11011000",	-- ##.##...
		2792 =>	"01101100",	-- .##.##..
		2793 =>	"00110110",	-- ..##.##.
		2794 =>	"00000000",	-- ........
		2795 =>	"00000000",	-- ........
		2796 =>	"00000000",	-- ........
		2797 =>	"00000000",	-- ........
		2798 =>	"00000000",	-- ........
		2799 =>	"00000000",	-- ........

		-- char 0xaf='\xaf
		2800 =>	"00000000",	-- ........
		2801 =>	"00000000",	-- ........
		2802 =>	"00000000",	-- ........
		2803 =>	"00000000",	-- ........
		2804 =>	"00000000",	-- ........
		2805 =>	"11011000",	-- ##.##...
		2806 =>	"01101100",	-- .##.##..
		2807 =>	"00110110",	-- ..##.##.
		2808 =>	"01101100",	-- .##.##..
		2809 =>	"11011000",	-- ##.##...
		2810 =>	"00000000",	-- ........
		2811 =>	"00000000",	-- ........
		2812 =>	"00000000",	-- ........
		2813 =>	"00000000",	-- ........
		2814 =>	"00000000",	-- ........
		2815 =>	"00000000",	-- ........

		-- char 0xb0='\xb0
		2816 =>	"01000100",	-- .#...#..
		2817 =>	"00010001",	-- ...#...#
		2818 =>	"01000100",	-- .#...#..
		2819 =>	"00010001",	-- ...#...#
		2820 =>	"01000100",	-- .#...#..
		2821 =>	"00010001",	-- ...#...#
		2822 =>	"01000100",	-- .#...#..
		2823 =>	"00010001",	-- ...#...#
		2824 =>	"01000100",	-- .#...#..
		2825 =>	"00010001",	-- ...#...#
		2826 =>	"01000100",	-- .#...#..
		2827 =>	"00010001",	-- ...#...#
		2828 =>	"01000100",	-- .#...#..
		2829 =>	"00010001",	-- ...#...#
		2830 =>	"01000100",	-- .#...#..
		2831 =>	"00010001",	-- ...#...#

		-- char 0xb1='\xb1
		2832 =>	"10101010",	-- #.#.#.#.
		2833 =>	"01010101",	-- .#.#.#.#
		2834 =>	"10101010",	-- #.#.#.#.
		2835 =>	"01010101",	-- .#.#.#.#
		2836 =>	"10101010",	-- #.#.#.#.
		2837 =>	"01010101",	-- .#.#.#.#
		2838 =>	"10101010",	-- #.#.#.#.
		2839 =>	"01010101",	-- .#.#.#.#
		2840 =>	"10101010",	-- #.#.#.#.
		2841 =>	"01010101",	-- .#.#.#.#
		2842 =>	"10101010",	-- #.#.#.#.
		2843 =>	"01010101",	-- .#.#.#.#
		2844 =>	"10101010",	-- #.#.#.#.
		2845 =>	"01010101",	-- .#.#.#.#
		2846 =>	"10101010",	-- #.#.#.#.
		2847 =>	"01010101",	-- .#.#.#.#

		-- char 0xb2='\xb2
		2848 =>	"01110111",	-- .###.###
		2849 =>	"11011101",	-- ##.###.#
		2850 =>	"01110111",	-- .###.###
		2851 =>	"11011101",	-- ##.###.#
		2852 =>	"01110111",	-- .###.###
		2853 =>	"11011101",	-- ##.###.#
		2854 =>	"01110111",	-- .###.###
		2855 =>	"11011101",	-- ##.###.#
		2856 =>	"01110111",	-- .###.###
		2857 =>	"11011101",	-- ##.###.#
		2858 =>	"01110111",	-- .###.###
		2859 =>	"11011101",	-- ##.###.#
		2860 =>	"01110111",	-- .###.###
		2861 =>	"11011101",	-- ##.###.#
		2862 =>	"01110111",	-- .###.###
		2863 =>	"11011101",	-- ##.###.#

		-- char 0xb3='\xb3
		2864 =>	"00011000",	-- ...##...
		2865 =>	"00011000",	-- ...##...
		2866 =>	"00011000",	-- ...##...
		2867 =>	"00011000",	-- ...##...
		2868 =>	"00011000",	-- ...##...
		2869 =>	"00011000",	-- ...##...
		2870 =>	"00011000",	-- ...##...
		2871 =>	"00011000",	-- ...##...
		2872 =>	"00011000",	-- ...##...
		2873 =>	"00011000",	-- ...##...
		2874 =>	"00011000",	-- ...##...
		2875 =>	"00011000",	-- ...##...
		2876 =>	"00011000",	-- ...##...
		2877 =>	"00011000",	-- ...##...
		2878 =>	"00011000",	-- ...##...
		2879 =>	"00011000",	-- ...##...

		-- char 0xb4='\xb4
		2880 =>	"00011000",	-- ...##...
		2881 =>	"00011000",	-- ...##...
		2882 =>	"00011000",	-- ...##...
		2883 =>	"00011000",	-- ...##...
		2884 =>	"00011000",	-- ...##...
		2885 =>	"00011000",	-- ...##...
		2886 =>	"00011000",	-- ...##...
		2887 =>	"00011000",	-- ...##...
		2888 =>	"11111000",	-- #####...
		2889 =>	"00011000",	-- ...##...
		2890 =>	"00011000",	-- ...##...
		2891 =>	"00011000",	-- ...##...
		2892 =>	"00011000",	-- ...##...
		2893 =>	"00011000",	-- ...##...
		2894 =>	"00011000",	-- ...##...
		2895 =>	"00011000",	-- ...##...

		-- char 0xb5='\xb5
		2896 =>	"00011000",	-- ...##...
		2897 =>	"00011000",	-- ...##...
		2898 =>	"00011000",	-- ...##...
		2899 =>	"00011000",	-- ...##...
		2900 =>	"00011000",	-- ...##...
		2901 =>	"00011000",	-- ...##...
		2902 =>	"11111000",	-- #####...
		2903 =>	"00011000",	-- ...##...
		2904 =>	"11111000",	-- #####...
		2905 =>	"00011000",	-- ...##...
		2906 =>	"00011000",	-- ...##...
		2907 =>	"00011000",	-- ...##...
		2908 =>	"00011000",	-- ...##...
		2909 =>	"00011000",	-- ...##...
		2910 =>	"00011000",	-- ...##...
		2911 =>	"00011000",	-- ...##...

		-- char 0xb6='\xb6
		2912 =>	"00110110",	-- ..##.##.
		2913 =>	"00110110",	-- ..##.##.
		2914 =>	"00110110",	-- ..##.##.
		2915 =>	"00110110",	-- ..##.##.
		2916 =>	"00110110",	-- ..##.##.
		2917 =>	"00110110",	-- ..##.##.
		2918 =>	"00110110",	-- ..##.##.
		2919 =>	"00110110",	-- ..##.##.
		2920 =>	"11110110",	-- ####.##.
		2921 =>	"00110110",	-- ..##.##.
		2922 =>	"00110110",	-- ..##.##.
		2923 =>	"00110110",	-- ..##.##.
		2924 =>	"00110110",	-- ..##.##.
		2925 =>	"00110110",	-- ..##.##.
		2926 =>	"00110110",	-- ..##.##.
		2927 =>	"00110110",	-- ..##.##.

		-- char 0xb7='\xb7
		2928 =>	"00000000",	-- ........
		2929 =>	"00000000",	-- ........
		2930 =>	"00000000",	-- ........
		2931 =>	"00000000",	-- ........
		2932 =>	"00000000",	-- ........
		2933 =>	"00000000",	-- ........
		2934 =>	"00000000",	-- ........
		2935 =>	"00000000",	-- ........
		2936 =>	"11111110",	-- #######.
		2937 =>	"00110110",	-- ..##.##.
		2938 =>	"00110110",	-- ..##.##.
		2939 =>	"00110110",	-- ..##.##.
		2940 =>	"00110110",	-- ..##.##.
		2941 =>	"00110110",	-- ..##.##.
		2942 =>	"00110110",	-- ..##.##.
		2943 =>	"00110110",	-- ..##.##.

		-- char 0xb8='\xb8
		2944 =>	"00000000",	-- ........
		2945 =>	"00000000",	-- ........
		2946 =>	"00000000",	-- ........
		2947 =>	"00000000",	-- ........
		2948 =>	"00000000",	-- ........
		2949 =>	"00000000",	-- ........
		2950 =>	"11111000",	-- #####...
		2951 =>	"00011000",	-- ...##...
		2952 =>	"11111000",	-- #####...
		2953 =>	"00011000",	-- ...##...
		2954 =>	"00011000",	-- ...##...
		2955 =>	"00011000",	-- ...##...
		2956 =>	"00011000",	-- ...##...
		2957 =>	"00011000",	-- ...##...
		2958 =>	"00011000",	-- ...##...
		2959 =>	"00011000",	-- ...##...

		-- char 0xb9='\xb9
		2960 =>	"00110110",	-- ..##.##.
		2961 =>	"00110110",	-- ..##.##.
		2962 =>	"00110110",	-- ..##.##.
		2963 =>	"00110110",	-- ..##.##.
		2964 =>	"00110110",	-- ..##.##.
		2965 =>	"00110110",	-- ..##.##.
		2966 =>	"11110110",	-- ####.##.
		2967 =>	"00000110",	-- .....##.
		2968 =>	"11110110",	-- ####.##.
		2969 =>	"00110110",	-- ..##.##.
		2970 =>	"00110110",	-- ..##.##.
		2971 =>	"00110110",	-- ..##.##.
		2972 =>	"00110110",	-- ..##.##.
		2973 =>	"00110110",	-- ..##.##.
		2974 =>	"00110110",	-- ..##.##.
		2975 =>	"00110110",	-- ..##.##.

		-- char 0xba='\xba
		2976 =>	"00110110",	-- ..##.##.
		2977 =>	"00110110",	-- ..##.##.
		2978 =>	"00110110",	-- ..##.##.
		2979 =>	"00110110",	-- ..##.##.
		2980 =>	"00110110",	-- ..##.##.
		2981 =>	"00110110",	-- ..##.##.
		2982 =>	"00110110",	-- ..##.##.
		2983 =>	"00110110",	-- ..##.##.
		2984 =>	"00110110",	-- ..##.##.
		2985 =>	"00110110",	-- ..##.##.
		2986 =>	"00110110",	-- ..##.##.
		2987 =>	"00110110",	-- ..##.##.
		2988 =>	"00110110",	-- ..##.##.
		2989 =>	"00110110",	-- ..##.##.
		2990 =>	"00110110",	-- ..##.##.
		2991 =>	"00110110",	-- ..##.##.

		-- char 0xbb='\xbb
		2992 =>	"00000000",	-- ........
		2993 =>	"00000000",	-- ........
		2994 =>	"00000000",	-- ........
		2995 =>	"00000000",	-- ........
		2996 =>	"00000000",	-- ........
		2997 =>	"00000000",	-- ........
		2998 =>	"11111110",	-- #######.
		2999 =>	"00000110",	-- .....##.
		3000 =>	"11110110",	-- ####.##.
		3001 =>	"00110110",	-- ..##.##.
		3002 =>	"00110110",	-- ..##.##.
		3003 =>	"00110110",	-- ..##.##.
		3004 =>	"00110110",	-- ..##.##.
		3005 =>	"00110110",	-- ..##.##.
		3006 =>	"00110110",	-- ..##.##.
		3007 =>	"00110110",	-- ..##.##.

		-- char 0xbc='\xbc
		3008 =>	"00110110",	-- ..##.##.
		3009 =>	"00110110",	-- ..##.##.
		3010 =>	"00110110",	-- ..##.##.
		3011 =>	"00110110",	-- ..##.##.
		3012 =>	"00110110",	-- ..##.##.
		3013 =>	"00110110",	-- ..##.##.
		3014 =>	"11110110",	-- ####.##.
		3015 =>	"00000110",	-- .....##.
		3016 =>	"11111110",	-- #######.
		3017 =>	"00000000",	-- ........
		3018 =>	"00000000",	-- ........
		3019 =>	"00000000",	-- ........
		3020 =>	"00000000",	-- ........
		3021 =>	"00000000",	-- ........
		3022 =>	"00000000",	-- ........
		3023 =>	"00000000",	-- ........

		-- char 0xbd='\xbd
		3024 =>	"00110110",	-- ..##.##.
		3025 =>	"00110110",	-- ..##.##.
		3026 =>	"00110110",	-- ..##.##.
		3027 =>	"00110110",	-- ..##.##.
		3028 =>	"00110110",	-- ..##.##.
		3029 =>	"00110110",	-- ..##.##.
		3030 =>	"00110110",	-- ..##.##.
		3031 =>	"00110110",	-- ..##.##.
		3032 =>	"11111110",	-- #######.
		3033 =>	"00000000",	-- ........
		3034 =>	"00000000",	-- ........
		3035 =>	"00000000",	-- ........
		3036 =>	"00000000",	-- ........
		3037 =>	"00000000",	-- ........
		3038 =>	"00000000",	-- ........
		3039 =>	"00000000",	-- ........

		-- char 0xbe='\xbe
		3040 =>	"00011000",	-- ...##...
		3041 =>	"00011000",	-- ...##...
		3042 =>	"00011000",	-- ...##...
		3043 =>	"00011000",	-- ...##...
		3044 =>	"00011000",	-- ...##...
		3045 =>	"00011000",	-- ...##...
		3046 =>	"11111000",	-- #####...
		3047 =>	"00011000",	-- ...##...
		3048 =>	"11111000",	-- #####...
		3049 =>	"00000000",	-- ........
		3050 =>	"00000000",	-- ........
		3051 =>	"00000000",	-- ........
		3052 =>	"00000000",	-- ........
		3053 =>	"00000000",	-- ........
		3054 =>	"00000000",	-- ........
		3055 =>	"00000000",	-- ........

		-- char 0xbf='\xbf
		3056 =>	"00000000",	-- ........
		3057 =>	"00000000",	-- ........
		3058 =>	"00000000",	-- ........
		3059 =>	"00000000",	-- ........
		3060 =>	"00000000",	-- ........
		3061 =>	"00000000",	-- ........
		3062 =>	"00000000",	-- ........
		3063 =>	"00000000",	-- ........
		3064 =>	"11111000",	-- #####...
		3065 =>	"00011000",	-- ...##...
		3066 =>	"00011000",	-- ...##...
		3067 =>	"00011000",	-- ...##...
		3068 =>	"00011000",	-- ...##...
		3069 =>	"00011000",	-- ...##...
		3070 =>	"00011000",	-- ...##...
		3071 =>	"00011000",	-- ...##...

		-- char 0xc0='\xc0
		3072 =>	"00011000",	-- ...##...
		3073 =>	"00011000",	-- ...##...
		3074 =>	"00011000",	-- ...##...
		3075 =>	"00011000",	-- ...##...
		3076 =>	"00011000",	-- ...##...
		3077 =>	"00011000",	-- ...##...
		3078 =>	"00011000",	-- ...##...
		3079 =>	"00011000",	-- ...##...
		3080 =>	"00011111",	-- ...#####
		3081 =>	"00000000",	-- ........
		3082 =>	"00000000",	-- ........
		3083 =>	"00000000",	-- ........
		3084 =>	"00000000",	-- ........
		3085 =>	"00000000",	-- ........
		3086 =>	"00000000",	-- ........
		3087 =>	"00000000",	-- ........

		-- char 0xc1='\xc1
		3088 =>	"00011000",	-- ...##...
		3089 =>	"00011000",	-- ...##...
		3090 =>	"00011000",	-- ...##...
		3091 =>	"00011000",	-- ...##...
		3092 =>	"00011000",	-- ...##...
		3093 =>	"00011000",	-- ...##...
		3094 =>	"00011000",	-- ...##...
		3095 =>	"00011000",	-- ...##...
		3096 =>	"11111111",	-- ########
		3097 =>	"00000000",	-- ........
		3098 =>	"00000000",	-- ........
		3099 =>	"00000000",	-- ........
		3100 =>	"00000000",	-- ........
		3101 =>	"00000000",	-- ........
		3102 =>	"00000000",	-- ........
		3103 =>	"00000000",	-- ........

		-- char 0xc2='\xc2
		3104 =>	"00000000",	-- ........
		3105 =>	"00000000",	-- ........
		3106 =>	"00000000",	-- ........
		3107 =>	"00000000",	-- ........
		3108 =>	"00000000",	-- ........
		3109 =>	"00000000",	-- ........
		3110 =>	"00000000",	-- ........
		3111 =>	"00000000",	-- ........
		3112 =>	"11111111",	-- ########
		3113 =>	"00011000",	-- ...##...
		3114 =>	"00011000",	-- ...##...
		3115 =>	"00011000",	-- ...##...
		3116 =>	"00011000",	-- ...##...
		3117 =>	"00011000",	-- ...##...
		3118 =>	"00011000",	-- ...##...
		3119 =>	"00011000",	-- ...##...

		-- char 0xc3='\xc3
		3120 =>	"00011000",	-- ...##...
		3121 =>	"00011000",	-- ...##...
		3122 =>	"00011000",	-- ...##...
		3123 =>	"00011000",	-- ...##...
		3124 =>	"00011000",	-- ...##...
		3125 =>	"00011000",	-- ...##...
		3126 =>	"00011000",	-- ...##...
		3127 =>	"00011000",	-- ...##...
		3128 =>	"00011111",	-- ...#####
		3129 =>	"00011000",	-- ...##...
		3130 =>	"00011000",	-- ...##...
		3131 =>	"00011000",	-- ...##...
		3132 =>	"00011000",	-- ...##...
		3133 =>	"00011000",	-- ...##...
		3134 =>	"00011000",	-- ...##...
		3135 =>	"00011000",	-- ...##...

		-- char 0xc4='\xc4
		3136 =>	"00000000",	-- ........
		3137 =>	"00000000",	-- ........
		3138 =>	"00000000",	-- ........
		3139 =>	"00000000",	-- ........
		3140 =>	"00000000",	-- ........
		3141 =>	"00000000",	-- ........
		3142 =>	"00000000",	-- ........
		3143 =>	"00000000",	-- ........
		3144 =>	"11111111",	-- ########
		3145 =>	"00000000",	-- ........
		3146 =>	"00000000",	-- ........
		3147 =>	"00000000",	-- ........
		3148 =>	"00000000",	-- ........
		3149 =>	"00000000",	-- ........
		3150 =>	"00000000",	-- ........
		3151 =>	"00000000",	-- ........

		-- char 0xc5='\xc5
		3152 =>	"00011000",	-- ...##...
		3153 =>	"00011000",	-- ...##...
		3154 =>	"00011000",	-- ...##...
		3155 =>	"00011000",	-- ...##...
		3156 =>	"00011000",	-- ...##...
		3157 =>	"00011000",	-- ...##...
		3158 =>	"00011000",	-- ...##...
		3159 =>	"00011000",	-- ...##...
		3160 =>	"11111111",	-- ########
		3161 =>	"00011000",	-- ...##...
		3162 =>	"00011000",	-- ...##...
		3163 =>	"00011000",	-- ...##...
		3164 =>	"00011000",	-- ...##...
		3165 =>	"00011000",	-- ...##...
		3166 =>	"00011000",	-- ...##...
		3167 =>	"00011000",	-- ...##...

		-- char 0xc6='\xc6
		3168 =>	"00011000",	-- ...##...
		3169 =>	"00011000",	-- ...##...
		3170 =>	"00011000",	-- ...##...
		3171 =>	"00011000",	-- ...##...
		3172 =>	"00011000",	-- ...##...
		3173 =>	"00011000",	-- ...##...
		3174 =>	"00011111",	-- ...#####
		3175 =>	"00011000",	-- ...##...
		3176 =>	"00011111",	-- ...#####
		3177 =>	"00011000",	-- ...##...
		3178 =>	"00011000",	-- ...##...
		3179 =>	"00011000",	-- ...##...
		3180 =>	"00011000",	-- ...##...
		3181 =>	"00011000",	-- ...##...
		3182 =>	"00011000",	-- ...##...
		3183 =>	"00011000",	-- ...##...

		-- char 0xc7='\xc7
		3184 =>	"00110110",	-- ..##.##.
		3185 =>	"00110110",	-- ..##.##.
		3186 =>	"00110110",	-- ..##.##.
		3187 =>	"00110110",	-- ..##.##.
		3188 =>	"00110110",	-- ..##.##.
		3189 =>	"00110110",	-- ..##.##.
		3190 =>	"00110110",	-- ..##.##.
		3191 =>	"00110110",	-- ..##.##.
		3192 =>	"00110111",	-- ..##.###
		3193 =>	"00110110",	-- ..##.##.
		3194 =>	"00110110",	-- ..##.##.
		3195 =>	"00110110",	-- ..##.##.
		3196 =>	"00110110",	-- ..##.##.
		3197 =>	"00110110",	-- ..##.##.
		3198 =>	"00110110",	-- ..##.##.
		3199 =>	"00110110",	-- ..##.##.

		-- char 0xc8='\xc8
		3200 =>	"00110110",	-- ..##.##.
		3201 =>	"00110110",	-- ..##.##.
		3202 =>	"00110110",	-- ..##.##.
		3203 =>	"00110110",	-- ..##.##.
		3204 =>	"00110110",	-- ..##.##.
		3205 =>	"00110110",	-- ..##.##.
		3206 =>	"00110111",	-- ..##.###
		3207 =>	"00110000",	-- ..##....
		3208 =>	"00111111",	-- ..######
		3209 =>	"00000000",	-- ........
		3210 =>	"00000000",	-- ........
		3211 =>	"00000000",	-- ........
		3212 =>	"00000000",	-- ........
		3213 =>	"00000000",	-- ........
		3214 =>	"00000000",	-- ........
		3215 =>	"00000000",	-- ........

		-- char 0xc9='\xc9
		3216 =>	"00000000",	-- ........
		3217 =>	"00000000",	-- ........
		3218 =>	"00000000",	-- ........
		3219 =>	"00000000",	-- ........
		3220 =>	"00000000",	-- ........
		3221 =>	"00000000",	-- ........
		3222 =>	"00111111",	-- ..######
		3223 =>	"00110000",	-- ..##....
		3224 =>	"00110111",	-- ..##.###
		3225 =>	"00110110",	-- ..##.##.
		3226 =>	"00110110",	-- ..##.##.
		3227 =>	"00110110",	-- ..##.##.
		3228 =>	"00110110",	-- ..##.##.
		3229 =>	"00110110",	-- ..##.##.
		3230 =>	"00110110",	-- ..##.##.
		3231 =>	"00110110",	-- ..##.##.

		-- char 0xca='\xca
		3232 =>	"00110110",	-- ..##.##.
		3233 =>	"00110110",	-- ..##.##.
		3234 =>	"00110110",	-- ..##.##.
		3235 =>	"00110110",	-- ..##.##.
		3236 =>	"00110110",	-- ..##.##.
		3237 =>	"00110110",	-- ..##.##.
		3238 =>	"11110111",	-- ####.###
		3239 =>	"00000000",	-- ........
		3240 =>	"11111111",	-- ########
		3241 =>	"00000000",	-- ........
		3242 =>	"00000000",	-- ........
		3243 =>	"00000000",	-- ........
		3244 =>	"00000000",	-- ........
		3245 =>	"00000000",	-- ........
		3246 =>	"00000000",	-- ........
		3247 =>	"00000000",	-- ........

		-- char 0xcb='\xcb
		3248 =>	"00000000",	-- ........
		3249 =>	"00000000",	-- ........
		3250 =>	"00000000",	-- ........
		3251 =>	"00000000",	-- ........
		3252 =>	"00000000",	-- ........
		3253 =>	"00000000",	-- ........
		3254 =>	"11111111",	-- ########
		3255 =>	"00000000",	-- ........
		3256 =>	"11110111",	-- ####.###
		3257 =>	"00110110",	-- ..##.##.
		3258 =>	"00110110",	-- ..##.##.
		3259 =>	"00110110",	-- ..##.##.
		3260 =>	"00110110",	-- ..##.##.
		3261 =>	"00110110",	-- ..##.##.
		3262 =>	"00110110",	-- ..##.##.
		3263 =>	"00110110",	-- ..##.##.

		-- char 0xcc='\xcc
		3264 =>	"00110110",	-- ..##.##.
		3265 =>	"00110110",	-- ..##.##.
		3266 =>	"00110110",	-- ..##.##.
		3267 =>	"00110110",	-- ..##.##.
		3268 =>	"00110110",	-- ..##.##.
		3269 =>	"00110110",	-- ..##.##.
		3270 =>	"00110111",	-- ..##.###
		3271 =>	"00110000",	-- ..##....
		3272 =>	"00110111",	-- ..##.###
		3273 =>	"00110110",	-- ..##.##.
		3274 =>	"00110110",	-- ..##.##.
		3275 =>	"00110110",	-- ..##.##.
		3276 =>	"00110110",	-- ..##.##.
		3277 =>	"00110110",	-- ..##.##.
		3278 =>	"00110110",	-- ..##.##.
		3279 =>	"00110110",	-- ..##.##.

		-- char 0xcd='\xcd
		3280 =>	"00000000",	-- ........
		3281 =>	"00000000",	-- ........
		3282 =>	"00000000",	-- ........
		3283 =>	"00000000",	-- ........
		3284 =>	"00000000",	-- ........
		3285 =>	"00000000",	-- ........
		3286 =>	"11111111",	-- ########
		3287 =>	"00000000",	-- ........
		3288 =>	"11111111",	-- ########
		3289 =>	"00000000",	-- ........
		3290 =>	"00000000",	-- ........
		3291 =>	"00000000",	-- ........
		3292 =>	"00000000",	-- ........
		3293 =>	"00000000",	-- ........
		3294 =>	"00000000",	-- ........
		3295 =>	"00000000",	-- ........

		-- char 0xce='\xce
		3296 =>	"00110110",	-- ..##.##.
		3297 =>	"00110110",	-- ..##.##.
		3298 =>	"00110110",	-- ..##.##.
		3299 =>	"00110110",	-- ..##.##.
		3300 =>	"00110110",	-- ..##.##.
		3301 =>	"00110110",	-- ..##.##.
		3302 =>	"11110111",	-- ####.###
		3303 =>	"00000000",	-- ........
		3304 =>	"11110111",	-- ####.###
		3305 =>	"00110110",	-- ..##.##.
		3306 =>	"00110110",	-- ..##.##.
		3307 =>	"00110110",	-- ..##.##.
		3308 =>	"00110110",	-- ..##.##.
		3309 =>	"00110110",	-- ..##.##.
		3310 =>	"00110110",	-- ..##.##.
		3311 =>	"00110110",	-- ..##.##.

		-- char 0xcf='\xcf
		3312 =>	"00011000",	-- ...##...
		3313 =>	"00011000",	-- ...##...
		3314 =>	"00011000",	-- ...##...
		3315 =>	"00011000",	-- ...##...
		3316 =>	"00011000",	-- ...##...
		3317 =>	"00011000",	-- ...##...
		3318 =>	"11111111",	-- ########
		3319 =>	"00000000",	-- ........
		3320 =>	"11111111",	-- ########
		3321 =>	"00000000",	-- ........
		3322 =>	"00000000",	-- ........
		3323 =>	"00000000",	-- ........
		3324 =>	"00000000",	-- ........
		3325 =>	"00000000",	-- ........
		3326 =>	"00000000",	-- ........
		3327 =>	"00000000",	-- ........

		-- char 0xd0='\xd0
		3328 =>	"00110110",	-- ..##.##.
		3329 =>	"00110110",	-- ..##.##.
		3330 =>	"00110110",	-- ..##.##.
		3331 =>	"00110110",	-- ..##.##.
		3332 =>	"00110110",	-- ..##.##.
		3333 =>	"00110110",	-- ..##.##.
		3334 =>	"00110110",	-- ..##.##.
		3335 =>	"00110110",	-- ..##.##.
		3336 =>	"11111111",	-- ########
		3337 =>	"00000000",	-- ........
		3338 =>	"00000000",	-- ........
		3339 =>	"00000000",	-- ........
		3340 =>	"00000000",	-- ........
		3341 =>	"00000000",	-- ........
		3342 =>	"00000000",	-- ........
		3343 =>	"00000000",	-- ........

		-- char 0xd1='\xd1
		3344 =>	"00000000",	-- ........
		3345 =>	"00000000",	-- ........
		3346 =>	"00000000",	-- ........
		3347 =>	"00000000",	-- ........
		3348 =>	"00000000",	-- ........
		3349 =>	"00000000",	-- ........
		3350 =>	"11111111",	-- ########
		3351 =>	"00000000",	-- ........
		3352 =>	"11111111",	-- ########
		3353 =>	"00011000",	-- ...##...
		3354 =>	"00011000",	-- ...##...
		3355 =>	"00011000",	-- ...##...
		3356 =>	"00011000",	-- ...##...
		3357 =>	"00011000",	-- ...##...
		3358 =>	"00011000",	-- ...##...
		3359 =>	"00011000",	-- ...##...

		-- char 0xd2='\xd2
		3360 =>	"00000000",	-- ........
		3361 =>	"00000000",	-- ........
		3362 =>	"00000000",	-- ........
		3363 =>	"00000000",	-- ........
		3364 =>	"00000000",	-- ........
		3365 =>	"00000000",	-- ........
		3366 =>	"00000000",	-- ........
		3367 =>	"00000000",	-- ........
		3368 =>	"11111111",	-- ########
		3369 =>	"00110110",	-- ..##.##.
		3370 =>	"00110110",	-- ..##.##.
		3371 =>	"00110110",	-- ..##.##.
		3372 =>	"00110110",	-- ..##.##.
		3373 =>	"00110110",	-- ..##.##.
		3374 =>	"00110110",	-- ..##.##.
		3375 =>	"00110110",	-- ..##.##.

		-- char 0xd3='\xd3
		3376 =>	"00110110",	-- ..##.##.
		3377 =>	"00110110",	-- ..##.##.
		3378 =>	"00110110",	-- ..##.##.
		3379 =>	"00110110",	-- ..##.##.
		3380 =>	"00110110",	-- ..##.##.
		3381 =>	"00110110",	-- ..##.##.
		3382 =>	"00110110",	-- ..##.##.
		3383 =>	"00110110",	-- ..##.##.
		3384 =>	"00111111",	-- ..######
		3385 =>	"00000000",	-- ........
		3386 =>	"00000000",	-- ........
		3387 =>	"00000000",	-- ........
		3388 =>	"00000000",	-- ........
		3389 =>	"00000000",	-- ........
		3390 =>	"00000000",	-- ........
		3391 =>	"00000000",	-- ........

		-- char 0xd4='\xd4
		3392 =>	"00011000",	-- ...##...
		3393 =>	"00011000",	-- ...##...
		3394 =>	"00011000",	-- ...##...
		3395 =>	"00011000",	-- ...##...
		3396 =>	"00011000",	-- ...##...
		3397 =>	"00011000",	-- ...##...
		3398 =>	"00011111",	-- ...#####
		3399 =>	"00011000",	-- ...##...
		3400 =>	"00011111",	-- ...#####
		3401 =>	"00000000",	-- ........
		3402 =>	"00000000",	-- ........
		3403 =>	"00000000",	-- ........
		3404 =>	"00000000",	-- ........
		3405 =>	"00000000",	-- ........
		3406 =>	"00000000",	-- ........
		3407 =>	"00000000",	-- ........

		-- char 0xd5='\xd5
		3408 =>	"00000000",	-- ........
		3409 =>	"00000000",	-- ........
		3410 =>	"00000000",	-- ........
		3411 =>	"00000000",	-- ........
		3412 =>	"00000000",	-- ........
		3413 =>	"00000000",	-- ........
		3414 =>	"00011111",	-- ...#####
		3415 =>	"00011000",	-- ...##...
		3416 =>	"00011111",	-- ...#####
		3417 =>	"00011000",	-- ...##...
		3418 =>	"00011000",	-- ...##...
		3419 =>	"00011000",	-- ...##...
		3420 =>	"00011000",	-- ...##...
		3421 =>	"00011000",	-- ...##...
		3422 =>	"00011000",	-- ...##...
		3423 =>	"00011000",	-- ...##...

		-- char 0xd6='\xd6
		3424 =>	"00000000",	-- ........
		3425 =>	"00000000",	-- ........
		3426 =>	"00000000",	-- ........
		3427 =>	"00000000",	-- ........
		3428 =>	"00000000",	-- ........
		3429 =>	"00000000",	-- ........
		3430 =>	"00000000",	-- ........
		3431 =>	"00000000",	-- ........
		3432 =>	"00111111",	-- ..######
		3433 =>	"00110110",	-- ..##.##.
		3434 =>	"00110110",	-- ..##.##.
		3435 =>	"00110110",	-- ..##.##.
		3436 =>	"00110110",	-- ..##.##.
		3437 =>	"00110110",	-- ..##.##.
		3438 =>	"00110110",	-- ..##.##.
		3439 =>	"00110110",	-- ..##.##.

		-- char 0xd7='\xd7
		3440 =>	"00110110",	-- ..##.##.
		3441 =>	"00110110",	-- ..##.##.
		3442 =>	"00110110",	-- ..##.##.
		3443 =>	"00110110",	-- ..##.##.
		3444 =>	"00110110",	-- ..##.##.
		3445 =>	"00110110",	-- ..##.##.
		3446 =>	"00110110",	-- ..##.##.
		3447 =>	"00110110",	-- ..##.##.
		3448 =>	"11111111",	-- ########
		3449 =>	"00110110",	-- ..##.##.
		3450 =>	"00110110",	-- ..##.##.
		3451 =>	"00110110",	-- ..##.##.
		3452 =>	"00110110",	-- ..##.##.
		3453 =>	"00110110",	-- ..##.##.
		3454 =>	"00110110",	-- ..##.##.
		3455 =>	"00110110",	-- ..##.##.

		-- char 0xd8='\xd8
		3456 =>	"00011000",	-- ...##...
		3457 =>	"00011000",	-- ...##...
		3458 =>	"00011000",	-- ...##...
		3459 =>	"00011000",	-- ...##...
		3460 =>	"00011000",	-- ...##...
		3461 =>	"00011000",	-- ...##...
		3462 =>	"11111111",	-- ########
		3463 =>	"00011000",	-- ...##...
		3464 =>	"11111111",	-- ########
		3465 =>	"00011000",	-- ...##...
		3466 =>	"00011000",	-- ...##...
		3467 =>	"00011000",	-- ...##...
		3468 =>	"00011000",	-- ...##...
		3469 =>	"00011000",	-- ...##...
		3470 =>	"00011000",	-- ...##...
		3471 =>	"00011000",	-- ...##...

		-- char 0xd9='\xd9
		3472 =>	"00011000",	-- ...##...
		3473 =>	"00011000",	-- ...##...
		3474 =>	"00011000",	-- ...##...
		3475 =>	"00011000",	-- ...##...
		3476 =>	"00011000",	-- ...##...
		3477 =>	"00011000",	-- ...##...
		3478 =>	"00011000",	-- ...##...
		3479 =>	"00011000",	-- ...##...
		3480 =>	"11111000",	-- #####...
		3481 =>	"00000000",	-- ........
		3482 =>	"00000000",	-- ........
		3483 =>	"00000000",	-- ........
		3484 =>	"00000000",	-- ........
		3485 =>	"00000000",	-- ........
		3486 =>	"00000000",	-- ........
		3487 =>	"00000000",	-- ........

		-- char 0xda='\xda
		3488 =>	"00000000",	-- ........
		3489 =>	"00000000",	-- ........
		3490 =>	"00000000",	-- ........
		3491 =>	"00000000",	-- ........
		3492 =>	"00000000",	-- ........
		3493 =>	"00000000",	-- ........
		3494 =>	"00000000",	-- ........
		3495 =>	"00000000",	-- ........
		3496 =>	"00011111",	-- ...#####
		3497 =>	"00011000",	-- ...##...
		3498 =>	"00011000",	-- ...##...
		3499 =>	"00011000",	-- ...##...
		3500 =>	"00011000",	-- ...##...
		3501 =>	"00011000",	-- ...##...
		3502 =>	"00011000",	-- ...##...
		3503 =>	"00011000",	-- ...##...

		-- char 0xdb='\xdb
		3504 =>	"11111111",	-- ########
		3505 =>	"11111111",	-- ########
		3506 =>	"11111111",	-- ########
		3507 =>	"11111111",	-- ########
		3508 =>	"11111111",	-- ########
		3509 =>	"11111111",	-- ########
		3510 =>	"11111111",	-- ########
		3511 =>	"11111111",	-- ########
		3512 =>	"11111111",	-- ########
		3513 =>	"11111111",	-- ########
		3514 =>	"11111111",	-- ########
		3515 =>	"11111111",	-- ########
		3516 =>	"11111111",	-- ########
		3517 =>	"11111111",	-- ########
		3518 =>	"11111111",	-- ########
		3519 =>	"11111111",	-- ########

		-- char 0xdc='\xdc
		3520 =>	"00000000",	-- ........
		3521 =>	"00000000",	-- ........
		3522 =>	"00000000",	-- ........
		3523 =>	"00000000",	-- ........
		3524 =>	"00000000",	-- ........
		3525 =>	"00000000",	-- ........
		3526 =>	"00000000",	-- ........
		3527 =>	"00000000",	-- ........
		3528 =>	"11111111",	-- ########
		3529 =>	"11111111",	-- ########
		3530 =>	"11111111",	-- ########
		3531 =>	"11111111",	-- ########
		3532 =>	"11111111",	-- ########
		3533 =>	"11111111",	-- ########
		3534 =>	"11111111",	-- ########
		3535 =>	"11111111",	-- ########

		-- char 0xdd='\xdd
		3536 =>	"11110000",	-- ####....
		3537 =>	"11110000",	-- ####....
		3538 =>	"11110000",	-- ####....
		3539 =>	"11110000",	-- ####....
		3540 =>	"11110000",	-- ####....
		3541 =>	"11110000",	-- ####....
		3542 =>	"11110000",	-- ####....
		3543 =>	"11110000",	-- ####....
		3544 =>	"11110000",	-- ####....
		3545 =>	"11110000",	-- ####....
		3546 =>	"11110000",	-- ####....
		3547 =>	"11110000",	-- ####....
		3548 =>	"11110000",	-- ####....
		3549 =>	"11110000",	-- ####....
		3550 =>	"11110000",	-- ####....
		3551 =>	"11110000",	-- ####....

		-- char 0xde='\xde
		3552 =>	"00001111",	-- ....####
		3553 =>	"00001111",	-- ....####
		3554 =>	"00001111",	-- ....####
		3555 =>	"00001111",	-- ....####
		3556 =>	"00001111",	-- ....####
		3557 =>	"00001111",	-- ....####
		3558 =>	"00001111",	-- ....####
		3559 =>	"00001111",	-- ....####
		3560 =>	"00001111",	-- ....####
		3561 =>	"00001111",	-- ....####
		3562 =>	"00001111",	-- ....####
		3563 =>	"00001111",	-- ....####
		3564 =>	"00001111",	-- ....####
		3565 =>	"00001111",	-- ....####
		3566 =>	"00001111",	-- ....####
		3567 =>	"00001111",	-- ....####

		-- char 0xdf='\xdf
		3568 =>	"11111111",	-- ########
		3569 =>	"11111111",	-- ########
		3570 =>	"11111111",	-- ########
		3571 =>	"11111111",	-- ########
		3572 =>	"11111111",	-- ########
		3573 =>	"11111111",	-- ########
		3574 =>	"11111111",	-- ########
		3575 =>	"11111111",	-- ########
		3576 =>	"00000000",	-- ........
		3577 =>	"00000000",	-- ........
		3578 =>	"00000000",	-- ........
		3579 =>	"00000000",	-- ........
		3580 =>	"00000000",	-- ........
		3581 =>	"00000000",	-- ........
		3582 =>	"00000000",	-- ........
		3583 =>	"00000000",	-- ........

		-- char 0xe0='\xe0
		3584 =>	"00000000",	-- ........
		3585 =>	"00000000",	-- ........
		3586 =>	"00000000",	-- ........
		3587 =>	"00000000",	-- ........
		3588 =>	"00000000",	-- ........
		3589 =>	"00000000",	-- ........
		3590 =>	"01110110",	-- .###.##.
		3591 =>	"11011100",	-- ##.###..
		3592 =>	"11011000",	-- ##.##...
		3593 =>	"11011000",	-- ##.##...
		3594 =>	"11011100",	-- ##.###..
		3595 =>	"01110110",	-- .###.##.
		3596 =>	"00000000",	-- ........
		3597 =>	"00000000",	-- ........
		3598 =>	"00000000",	-- ........
		3599 =>	"00000000",	-- ........

		-- char 0xe1='\xe1
		3600 =>	"00000000",	-- ........
		3601 =>	"00000000",	-- ........
		3602 =>	"00000000",	-- ........
		3603 =>	"00000000",	-- ........
		3604 =>	"00000000",	-- ........
		3605 =>	"01111100",	-- .#####..
		3606 =>	"11000110",	-- ##...##.
		3607 =>	"11111100",	-- ######..
		3608 =>	"11000110",	-- ##...##.
		3609 =>	"11000110",	-- ##...##.
		3610 =>	"11111100",	-- ######..
		3611 =>	"11000000",	-- ##......
		3612 =>	"11000000",	-- ##......
		3613 =>	"01000000",	-- .#......
		3614 =>	"00000000",	-- ........
		3615 =>	"00000000",	-- ........

		-- char 0xe2='\xe2
		3616 =>	"00000000",	-- ........
		3617 =>	"00000000",	-- ........
		3618 =>	"00000000",	-- ........
		3619 =>	"11111110",	-- #######.
		3620 =>	"11000110",	-- ##...##.
		3621 =>	"11000110",	-- ##...##.
		3622 =>	"11000000",	-- ##......
		3623 =>	"11000000",	-- ##......
		3624 =>	"11000000",	-- ##......
		3625 =>	"11000000",	-- ##......
		3626 =>	"11000000",	-- ##......
		3627 =>	"11000000",	-- ##......
		3628 =>	"00000000",	-- ........
		3629 =>	"00000000",	-- ........
		3630 =>	"00000000",	-- ........
		3631 =>	"00000000",	-- ........

		-- char 0xe3='\xe3
		3632 =>	"00000000",	-- ........
		3633 =>	"00000000",	-- ........
		3634 =>	"00000000",	-- ........
		3635 =>	"00000000",	-- ........
		3636 =>	"00000000",	-- ........
		3637 =>	"11111110",	-- #######.
		3638 =>	"01101100",	-- .##.##..
		3639 =>	"01101100",	-- .##.##..
		3640 =>	"01101100",	-- .##.##..
		3641 =>	"01101100",	-- .##.##..
		3642 =>	"01101100",	-- .##.##..
		3643 =>	"01101100",	-- .##.##..
		3644 =>	"00000000",	-- ........
		3645 =>	"00000000",	-- ........
		3646 =>	"00000000",	-- ........
		3647 =>	"00000000",	-- ........

		-- char 0xe4='\xe4
		3648 =>	"00000000",	-- ........
		3649 =>	"00000000",	-- ........
		3650 =>	"00000000",	-- ........
		3651 =>	"11111110",	-- #######.
		3652 =>	"11000110",	-- ##...##.
		3653 =>	"01100000",	-- .##.....
		3654 =>	"00110000",	-- ..##....
		3655 =>	"00011000",	-- ...##...
		3656 =>	"00110000",	-- ..##....
		3657 =>	"01100000",	-- .##.....
		3658 =>	"11000110",	-- ##...##.
		3659 =>	"11111110",	-- #######.
		3660 =>	"00000000",	-- ........
		3661 =>	"00000000",	-- ........
		3662 =>	"00000000",	-- ........
		3663 =>	"00000000",	-- ........

		-- char 0xe5='\xe5
		3664 =>	"00000000",	-- ........
		3665 =>	"00000000",	-- ........
		3666 =>	"00000000",	-- ........
		3667 =>	"00000000",	-- ........
		3668 =>	"00000000",	-- ........
		3669 =>	"00000000",	-- ........
		3670 =>	"01111110",	-- .######.
		3671 =>	"11011000",	-- ##.##...
		3672 =>	"11011000",	-- ##.##...
		3673 =>	"11011000",	-- ##.##...
		3674 =>	"11011000",	-- ##.##...
		3675 =>	"01110000",	-- .###....
		3676 =>	"00000000",	-- ........
		3677 =>	"00000000",	-- ........
		3678 =>	"00000000",	-- ........
		3679 =>	"00000000",	-- ........

		-- char 0xe6='\xe6
		3680 =>	"00000000",	-- ........
		3681 =>	"00000000",	-- ........
		3682 =>	"00000000",	-- ........
		3683 =>	"00000000",	-- ........
		3684 =>	"00000000",	-- ........
		3685 =>	"01100110",	-- .##..##.
		3686 =>	"01100110",	-- .##..##.
		3687 =>	"01100110",	-- .##..##.
		3688 =>	"01100110",	-- .##..##.
		3689 =>	"01111100",	-- .#####..
		3690 =>	"01100000",	-- .##.....
		3691 =>	"01100000",	-- .##.....
		3692 =>	"11000000",	-- ##......
		3693 =>	"00000000",	-- ........
		3694 =>	"00000000",	-- ........
		3695 =>	"00000000",	-- ........

		-- char 0xe7='\xe7
		3696 =>	"00000000",	-- ........
		3697 =>	"00000000",	-- ........
		3698 =>	"00000000",	-- ........
		3699 =>	"00000000",	-- ........
		3700 =>	"00000000",	-- ........
		3701 =>	"01110110",	-- .###.##.
		3702 =>	"11011100",	-- ##.###..
		3703 =>	"00011000",	-- ...##...
		3704 =>	"00011000",	-- ...##...
		3705 =>	"00011000",	-- ...##...
		3706 =>	"00011000",	-- ...##...
		3707 =>	"00011000",	-- ...##...
		3708 =>	"00000000",	-- ........
		3709 =>	"00000000",	-- ........
		3710 =>	"00000000",	-- ........
		3711 =>	"00000000",	-- ........

		-- char 0xe8='\xe8
		3712 =>	"00000000",	-- ........
		3713 =>	"00000000",	-- ........
		3714 =>	"00000000",	-- ........
		3715 =>	"01111110",	-- .######.
		3716 =>	"00011000",	-- ...##...
		3717 =>	"00111100",	-- ..####..
		3718 =>	"01100110",	-- .##..##.
		3719 =>	"01100110",	-- .##..##.
		3720 =>	"01100110",	-- .##..##.
		3721 =>	"00111100",	-- ..####..
		3722 =>	"00011000",	-- ...##...
		3723 =>	"01111110",	-- .######.
		3724 =>	"00000000",	-- ........
		3725 =>	"00000000",	-- ........
		3726 =>	"00000000",	-- ........
		3727 =>	"00000000",	-- ........

		-- char 0xe9='\xe9
		3728 =>	"00000000",	-- ........
		3729 =>	"00000000",	-- ........
		3730 =>	"00000000",	-- ........
		3731 =>	"00111000",	-- ..###...
		3732 =>	"01101100",	-- .##.##..
		3733 =>	"11000110",	-- ##...##.
		3734 =>	"11000110",	-- ##...##.
		3735 =>	"11111110",	-- #######.
		3736 =>	"11000110",	-- ##...##.
		3737 =>	"11000110",	-- ##...##.
		3738 =>	"01101100",	-- .##.##..
		3739 =>	"00111000",	-- ..###...
		3740 =>	"00000000",	-- ........
		3741 =>	"00000000",	-- ........
		3742 =>	"00000000",	-- ........
		3743 =>	"00000000",	-- ........

		-- char 0xea='\xea
		3744 =>	"00000000",	-- ........
		3745 =>	"00000000",	-- ........
		3746 =>	"00000000",	-- ........
		3747 =>	"00111000",	-- ..###...
		3748 =>	"01101100",	-- .##.##..
		3749 =>	"11000110",	-- ##...##.
		3750 =>	"11000110",	-- ##...##.
		3751 =>	"11000110",	-- ##...##.
		3752 =>	"01101100",	-- .##.##..
		3753 =>	"01101100",	-- .##.##..
		3754 =>	"01101100",	-- .##.##..
		3755 =>	"11101110",	-- ###.###.
		3756 =>	"00000000",	-- ........
		3757 =>	"00000000",	-- ........
		3758 =>	"00000000",	-- ........
		3759 =>	"00000000",	-- ........

		-- char 0xeb='\xeb
		3760 =>	"00000000",	-- ........
		3761 =>	"00000000",	-- ........
		3762 =>	"00000000",	-- ........
		3763 =>	"00011110",	-- ...####.
		3764 =>	"00110000",	-- ..##....
		3765 =>	"00011000",	-- ...##...
		3766 =>	"00001100",	-- ....##..
		3767 =>	"00111110",	-- ..#####.
		3768 =>	"01100110",	-- .##..##.
		3769 =>	"01100110",	-- .##..##.
		3770 =>	"01100110",	-- .##..##.
		3771 =>	"00111100",	-- ..####..
		3772 =>	"00000000",	-- ........
		3773 =>	"00000000",	-- ........
		3774 =>	"00000000",	-- ........
		3775 =>	"00000000",	-- ........

		-- char 0xec='\xec
		3776 =>	"00000000",	-- ........
		3777 =>	"00000000",	-- ........
		3778 =>	"00000000",	-- ........
		3779 =>	"00000000",	-- ........
		3780 =>	"00000000",	-- ........
		3781 =>	"00000000",	-- ........
		3782 =>	"01111110",	-- .######.
		3783 =>	"11011011",	-- ##.##.##
		3784 =>	"11011011",	-- ##.##.##
		3785 =>	"01111110",	-- .######.
		3786 =>	"00000000",	-- ........
		3787 =>	"00000000",	-- ........
		3788 =>	"00000000",	-- ........
		3789 =>	"00000000",	-- ........
		3790 =>	"00000000",	-- ........
		3791 =>	"00000000",	-- ........

		-- char 0xed='\xed
		3792 =>	"00000000",	-- ........
		3793 =>	"00000000",	-- ........
		3794 =>	"00000000",	-- ........
		3795 =>	"00000011",	-- ......##
		3796 =>	"00000110",	-- .....##.
		3797 =>	"01111110",	-- .######.
		3798 =>	"11011011",	-- ##.##.##
		3799 =>	"11011011",	-- ##.##.##
		3800 =>	"11110011",	-- ####..##
		3801 =>	"01111110",	-- .######.
		3802 =>	"01100000",	-- .##.....
		3803 =>	"11000000",	-- ##......
		3804 =>	"00000000",	-- ........
		3805 =>	"00000000",	-- ........
		3806 =>	"00000000",	-- ........
		3807 =>	"00000000",	-- ........

		-- char 0xee='\xee
		3808 =>	"00000000",	-- ........
		3809 =>	"00000000",	-- ........
		3810 =>	"00000000",	-- ........
		3811 =>	"00011100",	-- ...###..
		3812 =>	"00110000",	-- ..##....
		3813 =>	"01100000",	-- .##.....
		3814 =>	"01100000",	-- .##.....
		3815 =>	"01111100",	-- .#####..
		3816 =>	"01100000",	-- .##.....
		3817 =>	"01100000",	-- .##.....
		3818 =>	"00110000",	-- ..##....
		3819 =>	"00011100",	-- ...###..
		3820 =>	"00000000",	-- ........
		3821 =>	"00000000",	-- ........
		3822 =>	"00000000",	-- ........
		3823 =>	"00000000",	-- ........

		-- char 0xef='\xef
		3824 =>	"00000000",	-- ........
		3825 =>	"00000000",	-- ........
		3826 =>	"00000000",	-- ........
		3827 =>	"00000000",	-- ........
		3828 =>	"01111100",	-- .#####..
		3829 =>	"11000110",	-- ##...##.
		3830 =>	"11000110",	-- ##...##.
		3831 =>	"11000110",	-- ##...##.
		3832 =>	"11000110",	-- ##...##.
		3833 =>	"11000110",	-- ##...##.
		3834 =>	"11000110",	-- ##...##.
		3835 =>	"11000110",	-- ##...##.
		3836 =>	"00000000",	-- ........
		3837 =>	"00000000",	-- ........
		3838 =>	"00000000",	-- ........
		3839 =>	"00000000",	-- ........

		-- char 0xf0='\xf0
		3840 =>	"00000000",	-- ........
		3841 =>	"00000000",	-- ........
		3842 =>	"00000000",	-- ........
		3843 =>	"00000000",	-- ........
		3844 =>	"11111110",	-- #######.
		3845 =>	"00000000",	-- ........
		3846 =>	"00000000",	-- ........
		3847 =>	"11111110",	-- #######.
		3848 =>	"00000000",	-- ........
		3849 =>	"00000000",	-- ........
		3850 =>	"11111110",	-- #######.
		3851 =>	"00000000",	-- ........
		3852 =>	"00000000",	-- ........
		3853 =>	"00000000",	-- ........
		3854 =>	"00000000",	-- ........
		3855 =>	"00000000",	-- ........

		-- char 0xf1='\xf1
		3856 =>	"00000000",	-- ........
		3857 =>	"00000000",	-- ........
		3858 =>	"00000000",	-- ........
		3859 =>	"00000000",	-- ........
		3860 =>	"00011000",	-- ...##...
		3861 =>	"00011000",	-- ...##...
		3862 =>	"01111110",	-- .######.
		3863 =>	"00011000",	-- ...##...
		3864 =>	"00011000",	-- ...##...
		3865 =>	"00000000",	-- ........
		3866 =>	"00000000",	-- ........
		3867 =>	"11111111",	-- ########
		3868 =>	"00000000",	-- ........
		3869 =>	"00000000",	-- ........
		3870 =>	"00000000",	-- ........
		3871 =>	"00000000",	-- ........

		-- char 0xf2='\xf2
		3872 =>	"00000000",	-- ........
		3873 =>	"00000000",	-- ........
		3874 =>	"00000000",	-- ........
		3875 =>	"00110000",	-- ..##....
		3876 =>	"00011000",	-- ...##...
		3877 =>	"00001100",	-- ....##..
		3878 =>	"00000110",	-- .....##.
		3879 =>	"00001100",	-- ....##..
		3880 =>	"00011000",	-- ...##...
		3881 =>	"00110000",	-- ..##....
		3882 =>	"00000000",	-- ........
		3883 =>	"01111110",	-- .######.
		3884 =>	"00000000",	-- ........
		3885 =>	"00000000",	-- ........
		3886 =>	"00000000",	-- ........
		3887 =>	"00000000",	-- ........

		-- char 0xf3='\xf3
		3888 =>	"00000000",	-- ........
		3889 =>	"00000000",	-- ........
		3890 =>	"00000000",	-- ........
		3891 =>	"00001100",	-- ....##..
		3892 =>	"00011000",	-- ...##...
		3893 =>	"00110000",	-- ..##....
		3894 =>	"01100000",	-- .##.....
		3895 =>	"00110000",	-- ..##....
		3896 =>	"00011000",	-- ...##...
		3897 =>	"00001100",	-- ....##..
		3898 =>	"00000000",	-- ........
		3899 =>	"01111110",	-- .######.
		3900 =>	"00000000",	-- ........
		3901 =>	"00000000",	-- ........
		3902 =>	"00000000",	-- ........
		3903 =>	"00000000",	-- ........

		-- char 0xf4='\xf4
		3904 =>	"00000000",	-- ........
		3905 =>	"00000000",	-- ........
		3906 =>	"00000000",	-- ........
		3907 =>	"00001110",	-- ....###.
		3908 =>	"00011011",	-- ...##.##
		3909 =>	"00011011",	-- ...##.##
		3910 =>	"00011000",	-- ...##...
		3911 =>	"00011000",	-- ...##...
		3912 =>	"00011000",	-- ...##...
		3913 =>	"00011000",	-- ...##...
		3914 =>	"00011000",	-- ...##...
		3915 =>	"00011000",	-- ...##...
		3916 =>	"00011000",	-- ...##...
		3917 =>	"00011000",	-- ...##...
		3918 =>	"00011000",	-- ...##...
		3919 =>	"00011000",	-- ...##...

		-- char 0xf5='\xf5
		3920 =>	"00011000",	-- ...##...
		3921 =>	"00011000",	-- ...##...
		3922 =>	"00011000",	-- ...##...
		3923 =>	"00011000",	-- ...##...
		3924 =>	"00011000",	-- ...##...
		3925 =>	"00011000",	-- ...##...
		3926 =>	"00011000",	-- ...##...
		3927 =>	"00011000",	-- ...##...
		3928 =>	"00011000",	-- ...##...
		3929 =>	"11011000",	-- ##.##...
		3930 =>	"11011000",	-- ##.##...
		3931 =>	"01110000",	-- .###....
		3932 =>	"00000000",	-- ........
		3933 =>	"00000000",	-- ........
		3934 =>	"00000000",	-- ........
		3935 =>	"00000000",	-- ........

		-- char 0xf6='\xf6
		3936 =>	"00000000",	-- ........
		3937 =>	"00000000",	-- ........
		3938 =>	"00000000",	-- ........
		3939 =>	"00000000",	-- ........
		3940 =>	"00011000",	-- ...##...
		3941 =>	"00011000",	-- ...##...
		3942 =>	"00000000",	-- ........
		3943 =>	"01111110",	-- .######.
		3944 =>	"00000000",	-- ........
		3945 =>	"00011000",	-- ...##...
		3946 =>	"00011000",	-- ...##...
		3947 =>	"00000000",	-- ........
		3948 =>	"00000000",	-- ........
		3949 =>	"00000000",	-- ........
		3950 =>	"00000000",	-- ........
		3951 =>	"00000000",	-- ........

		-- char 0xf7='\xf7
		3952 =>	"00000000",	-- ........
		3953 =>	"00000000",	-- ........
		3954 =>	"00000000",	-- ........
		3955 =>	"00000000",	-- ........
		3956 =>	"00000000",	-- ........
		3957 =>	"01110110",	-- .###.##.
		3958 =>	"11011100",	-- ##.###..
		3959 =>	"00000000",	-- ........
		3960 =>	"01110110",	-- .###.##.
		3961 =>	"11011100",	-- ##.###..
		3962 =>	"00000000",	-- ........
		3963 =>	"00000000",	-- ........
		3964 =>	"00000000",	-- ........
		3965 =>	"00000000",	-- ........
		3966 =>	"00000000",	-- ........
		3967 =>	"00000000",	-- ........

		-- char 0xf8='\xf8
		3968 =>	"00000000",	-- ........
		3969 =>	"00000000",	-- ........
		3970 =>	"00111000",	-- ..###...
		3971 =>	"01101100",	-- .##.##..
		3972 =>	"01101100",	-- .##.##..
		3973 =>	"00111000",	-- ..###...
		3974 =>	"00000000",	-- ........
		3975 =>	"00000000",	-- ........
		3976 =>	"00000000",	-- ........
		3977 =>	"00000000",	-- ........
		3978 =>	"00000000",	-- ........
		3979 =>	"00000000",	-- ........
		3980 =>	"00000000",	-- ........
		3981 =>	"00000000",	-- ........
		3982 =>	"00000000",	-- ........
		3983 =>	"00000000",	-- ........

		-- char 0xf9='\xf9
		3984 =>	"00000000",	-- ........
		3985 =>	"00000000",	-- ........
		3986 =>	"00000000",	-- ........
		3987 =>	"00000000",	-- ........
		3988 =>	"00000000",	-- ........
		3989 =>	"00000000",	-- ........
		3990 =>	"00000000",	-- ........
		3991 =>	"00011000",	-- ...##...
		3992 =>	"00011000",	-- ...##...
		3993 =>	"00000000",	-- ........
		3994 =>	"00000000",	-- ........
		3995 =>	"00000000",	-- ........
		3996 =>	"00000000",	-- ........
		3997 =>	"00000000",	-- ........
		3998 =>	"00000000",	-- ........
		3999 =>	"00000000",	-- ........

		-- char 0xfa='\xfa
		4000 =>	"00000000",	-- ........
		4001 =>	"00000000",	-- ........
		4002 =>	"00000000",	-- ........
		4003 =>	"00000000",	-- ........
		4004 =>	"00000000",	-- ........
		4005 =>	"00000000",	-- ........
		4006 =>	"00000000",	-- ........
		4007 =>	"00000000",	-- ........
		4008 =>	"00011000",	-- ...##...
		4009 =>	"00000000",	-- ........
		4010 =>	"00000000",	-- ........
		4011 =>	"00000000",	-- ........
		4012 =>	"00000000",	-- ........
		4013 =>	"00000000",	-- ........
		4014 =>	"00000000",	-- ........
		4015 =>	"00000000",	-- ........

		-- char 0xfb='\xfb
		4016 =>	"00000000",	-- ........
		4017 =>	"00000000",	-- ........
		4018 =>	"00001111",	-- ....####
		4019 =>	"00001100",	-- ....##..
		4020 =>	"00001100",	-- ....##..
		4021 =>	"00001100",	-- ....##..
		4022 =>	"00001100",	-- ....##..
		4023 =>	"00001100",	-- ....##..
		4024 =>	"11101100",	-- ###.##..
		4025 =>	"01101100",	-- .##.##..
		4026 =>	"00111100",	-- ..####..
		4027 =>	"00011100",	-- ...###..
		4028 =>	"00000000",	-- ........
		4029 =>	"00000000",	-- ........
		4030 =>	"00000000",	-- ........
		4031 =>	"00000000",	-- ........

		-- char 0xfc='\xfc
		4032 =>	"00000000",	-- ........
		4033 =>	"00000000",	-- ........
		4034 =>	"11011000",	-- ##.##...
		4035 =>	"01101100",	-- .##.##..
		4036 =>	"01101100",	-- .##.##..
		4037 =>	"01101100",	-- .##.##..
		4038 =>	"01101100",	-- .##.##..
		4039 =>	"01101100",	-- .##.##..
		4040 =>	"00000000",	-- ........
		4041 =>	"00000000",	-- ........
		4042 =>	"00000000",	-- ........
		4043 =>	"00000000",	-- ........
		4044 =>	"00000000",	-- ........
		4045 =>	"00000000",	-- ........
		4046 =>	"00000000",	-- ........
		4047 =>	"00000000",	-- ........

		-- char 0xfd='\xfd
		4048 =>	"00000000",	-- ........
		4049 =>	"00000000",	-- ........
		4050 =>	"01110000",	-- .###....
		4051 =>	"11011000",	-- ##.##...
		4052 =>	"00110000",	-- ..##....
		4053 =>	"01100000",	-- .##.....
		4054 =>	"11001000",	-- ##..#...
		4055 =>	"11111000",	-- #####...
		4056 =>	"00000000",	-- ........
		4057 =>	"00000000",	-- ........
		4058 =>	"00000000",	-- ........
		4059 =>	"00000000",	-- ........
		4060 =>	"00000000",	-- ........
		4061 =>	"00000000",	-- ........
		4062 =>	"00000000",	-- ........
		4063 =>	"00000000",	-- ........

		-- char 0xfe='\xfe
		4064 =>	"00000000",	-- ........
		4065 =>	"00000000",	-- ........
		4066 =>	"00000000",	-- ........
		4067 =>	"00000000",	-- ........
		4068 =>	"00000000",	-- ........
		4069 =>	"01111100",	-- .#####..
		4070 =>	"01111100",	-- .#####..
		4071 =>	"01111100",	-- .#####..
		4072 =>	"01111100",	-- .#####..
		4073 =>	"01111100",	-- .#####..
		4074 =>	"01111100",	-- .#####..
		4075 =>	"00000000",	-- ........
		4076 =>	"00000000",	-- ........
		4077 =>	"00000000",	-- ........
		4078 =>	"00000000",	-- ........
		4079 =>	"00000000",	-- ........

		-- char 0xff='\xff
		4080 =>	"00000000",	-- ........
		4081 =>	"00000000",	-- ........
		4082 =>	"00000000",	-- ........
		4083 =>	"00000000",	-- ........
		4084 =>	"00000000",	-- ........
		4085 =>	"00000000",	-- ........
		4086 =>	"00000000",	-- ........
		4087 =>	"00000000",	-- ........
		4088 =>	"00000000",	-- ........
		4089 =>	"00000000",	-- ........
		4090 =>	"00000000",	-- ........
		4091 =>	"00000000",	-- ........
		4092 =>	"00000000",	-- ........
		4093 =>	"00000000",	-- ........
		4094 =>	"00000000",	-- ........
		4095 =>	"00000000",	-- ........
	others => (others => '0')
    );

end font8x16_xark;
