library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.font_block_pack.all;

package font8x8_xark is

constant font8x8_block : font8_block_type := (
		-- char 0x00='\0' 
		0 =>	"00000000",	-- ........
		1 =>	"00000000",	-- ........
		2 =>	"00000000",	-- ........
		3 =>	"00000000",	-- ........
		4 =>	"00000000",	-- ........
		5 =>	"00000000",	-- ........
		6 =>	"00000000",	-- ........
		7 =>	"00000000",	-- ........

		-- char 0x01='\x01
		8 =>	"01111110",	-- .######.
		9 =>	"10000001",	-- #......#
		10 =>	"10100101",	-- #.#..#.#
		11 =>	"10000001",	-- #......#
		12 =>	"10111101",	-- #.####.#
		13 =>	"10011001",	-- #..##..#
		14 =>	"10000001",	-- #......#
		15 =>	"01111110",	-- .######.

		-- char 0x02='\x02
		16 =>	"01111110",	-- .######.
		17 =>	"11111111",	-- ########
		18 =>	"11011011",	-- ##.##.##
		19 =>	"11111111",	-- ########
		20 =>	"11000011",	-- ##....##
		21 =>	"11100111",	-- ###..###
		22 =>	"11111111",	-- ########
		23 =>	"01111110",	-- .######.

		-- char 0x03='\x03
		24 =>	"01101100",	-- .##.##..
		25 =>	"11111110",	-- #######.
		26 =>	"11111110",	-- #######.
		27 =>	"11111110",	-- #######.
		28 =>	"01111100",	-- .#####..
		29 =>	"00111000",	-- ..###...
		30 =>	"00010000",	-- ...#....
		31 =>	"00000000",	-- ........

		-- char 0x04='\x04
		32 =>	"00010000",	-- ...#....
		33 =>	"00111000",	-- ..###...
		34 =>	"01111100",	-- .#####..
		35 =>	"11111110",	-- #######.
		36 =>	"01111100",	-- .#####..
		37 =>	"00111000",	-- ..###...
		38 =>	"00010000",	-- ...#....
		39 =>	"00000000",	-- ........

		-- char 0x05='\x05
		40 =>	"00111000",	-- ..###...
		41 =>	"01111100",	-- .#####..
		42 =>	"00111000",	-- ..###...
		43 =>	"11111110",	-- #######.
		44 =>	"11111110",	-- #######.
		45 =>	"11010110",	-- ##.#.##.
		46 =>	"00010000",	-- ...#....
		47 =>	"00111000",	-- ..###...

		-- char 0x06='\x06
		48 =>	"00010000",	-- ...#....
		49 =>	"00111000",	-- ..###...
		50 =>	"01111100",	-- .#####..
		51 =>	"11111110",	-- #######.
		52 =>	"11111110",	-- #######.
		53 =>	"01010100",	-- .#.#.#..
		54 =>	"00010000",	-- ...#....
		55 =>	"00111000",	-- ..###...

		-- char 0x07='\a' 
		56 =>	"00000000",	-- ........
		57 =>	"00000000",	-- ........
		58 =>	"00011000",	-- ...##...
		59 =>	"00111100",	-- ..####..
		60 =>	"00111100",	-- ..####..
		61 =>	"00011000",	-- ...##...
		62 =>	"00000000",	-- ........
		63 =>	"00000000",	-- ........

		-- char 0x08='\b' 
		64 =>	"11111111",	-- ########
		65 =>	"11111111",	-- ########
		66 =>	"11100111",	-- ###..###
		67 =>	"11000011",	-- ##....##
		68 =>	"11000011",	-- ##....##
		69 =>	"11100111",	-- ###..###
		70 =>	"11111111",	-- ########
		71 =>	"11111111",	-- ########

		-- char 0x09='\t' 
		72 =>	"00000000",	-- ........
		73 =>	"00111100",	-- ..####..
		74 =>	"01100110",	-- .##..##.
		75 =>	"01000010",	-- .#....#.
		76 =>	"01000010",	-- .#....#.
		77 =>	"01100110",	-- .##..##.
		78 =>	"00111100",	-- ..####..
		79 =>	"00000000",	-- ........

		-- char 0x0a='\n' 
		80 =>	"11111111",	-- ########
		81 =>	"11000011",	-- ##....##
		82 =>	"10011001",	-- #..##..#
		83 =>	"10111101",	-- #.####.#
		84 =>	"10111101",	-- #.####.#
		85 =>	"10011001",	-- #..##..#
		86 =>	"11000011",	-- ##....##
		87 =>	"11111111",	-- ########

		-- char 0x0b='\v' 
		88 =>	"00001111",	-- ....####
		89 =>	"00000111",	-- .....###
		90 =>	"00001111",	-- ....####
		91 =>	"01111101",	-- .#####.#
		92 =>	"11001100",	-- ##..##..
		93 =>	"11001100",	-- ##..##..
		94 =>	"11001100",	-- ##..##..
		95 =>	"01111000",	-- .####...

		-- char 0x0c='\f' 
		96 =>	"00111100",	-- ..####..
		97 =>	"01100110",	-- .##..##.
		98 =>	"01100110",	-- .##..##.
		99 =>	"01100110",	-- .##..##.
		100 =>	"00111100",	-- ..####..
		101 =>	"00011000",	-- ...##...
		102 =>	"01111110",	-- .######.
		103 =>	"00011000",	-- ...##...

		-- char 0x0d='\r' 
		104 =>	"00111111",	-- ..######
		105 =>	"00110011",	-- ..##..##
		106 =>	"00111111",	-- ..######
		107 =>	"00110000",	-- ..##....
		108 =>	"00110000",	-- ..##....
		109 =>	"01110000",	-- .###....
		110 =>	"11110000",	-- ####....
		111 =>	"11100000",	-- ###.....

		-- char 0x0e='\x0e
		112 =>	"01111111",	-- .#######
		113 =>	"01100011",	-- .##...##
		114 =>	"01111111",	-- .#######
		115 =>	"01100011",	-- .##...##
		116 =>	"01100011",	-- .##...##
		117 =>	"01100111",	-- .##..###
		118 =>	"11100110",	-- ###..##.
		119 =>	"11000000",	-- ##......

		-- char 0x0f='\x0f
		120 =>	"10011001",	-- #..##..#
		121 =>	"01011010",	-- .#.##.#.
		122 =>	"00111100",	-- ..####..
		123 =>	"11100111",	-- ###..###
		124 =>	"11100111",	-- ###..###
		125 =>	"00111100",	-- ..####..
		126 =>	"01011010",	-- .#.##.#.
		127 =>	"10011001",	-- #..##..#

		-- char 0x10='\x10
		128 =>	"11000000",	-- ##......
		129 =>	"11110000",	-- ####....
		130 =>	"11111100",	-- ######..
		131 =>	"11111111",	-- ########
		132 =>	"11111111",	-- ########
		133 =>	"11111100",	-- ######..
		134 =>	"11110000",	-- ####....
		135 =>	"11000000",	-- ##......

		-- char 0x11='\x11
		136 =>	"00000011",	-- ......##
		137 =>	"00001111",	-- ....####
		138 =>	"00111111",	-- ..######
		139 =>	"11111111",	-- ########
		140 =>	"11111111",	-- ########
		141 =>	"00111111",	-- ..######
		142 =>	"00001111",	-- ....####
		143 =>	"00000011",	-- ......##

		-- char 0x12='\x12
		144 =>	"00011000",	-- ...##...
		145 =>	"00111100",	-- ..####..
		146 =>	"01111110",	-- .######.
		147 =>	"00011000",	-- ...##...
		148 =>	"00011000",	-- ...##...
		149 =>	"01111110",	-- .######.
		150 =>	"00111100",	-- ..####..
		151 =>	"00011000",	-- ...##...

		-- char 0x13='\x13
		152 =>	"01100110",	-- .##..##.
		153 =>	"01100110",	-- .##..##.
		154 =>	"01100110",	-- .##..##.
		155 =>	"01100110",	-- .##..##.
		156 =>	"01100110",	-- .##..##.
		157 =>	"00000000",	-- ........
		158 =>	"01100110",	-- .##..##.
		159 =>	"00000000",	-- ........

		-- char 0x14='\x14
		160 =>	"01111111",	-- .#######
		161 =>	"11011011",	-- ##.##.##
		162 =>	"11011011",	-- ##.##.##
		163 =>	"01111011",	-- .####.##
		164 =>	"00011011",	-- ...##.##
		165 =>	"00011011",	-- ...##.##
		166 =>	"00011011",	-- ...##.##
		167 =>	"00000000",	-- ........

		-- char 0x15='\x15
		168 =>	"01111110",	-- .######.
		169 =>	"11000011",	-- ##....##
		170 =>	"01111000",	-- .####...
		171 =>	"11001100",	-- ##..##..
		172 =>	"11001100",	-- ##..##..
		173 =>	"01111000",	-- .####...
		174 =>	"10001100",	-- #...##..
		175 =>	"11111000",	-- #####...

		-- char 0x16='\x16
		176 =>	"00000000",	-- ........
		177 =>	"00000000",	-- ........
		178 =>	"00000000",	-- ........
		179 =>	"00000000",	-- ........
		180 =>	"01111110",	-- .######.
		181 =>	"01111110",	-- .######.
		182 =>	"01111110",	-- .######.
		183 =>	"00000000",	-- ........

		-- char 0x17='\x17
		184 =>	"00011000",	-- ...##...
		185 =>	"00111100",	-- ..####..
		186 =>	"01111110",	-- .######.
		187 =>	"00011000",	-- ...##...
		188 =>	"01111110",	-- .######.
		189 =>	"00111100",	-- ..####..
		190 =>	"00011000",	-- ...##...
		191 =>	"11111111",	-- ########

		-- char 0x18='\x18
		192 =>	"00011000",	-- ...##...
		193 =>	"00111100",	-- ..####..
		194 =>	"01111110",	-- .######.
		195 =>	"00011000",	-- ...##...
		196 =>	"00011000",	-- ...##...
		197 =>	"00011000",	-- ...##...
		198 =>	"00011000",	-- ...##...
		199 =>	"00011000",	-- ...##...

		-- char 0x19='\x19
		200 =>	"00011000",	-- ...##...
		201 =>	"00011000",	-- ...##...
		202 =>	"00011000",	-- ...##...
		203 =>	"00011000",	-- ...##...
		204 =>	"00011000",	-- ...##...
		205 =>	"01111110",	-- .######.
		206 =>	"00111100",	-- ..####..
		207 =>	"00011000",	-- ...##...

		-- char 0x1a='\x1a
		208 =>	"00000000",	-- ........
		209 =>	"00000100",	-- .....#..
		210 =>	"00000110",	-- .....##.
		211 =>	"11111111",	-- ########
		212 =>	"11111111",	-- ########
		213 =>	"00000110",	-- .....##.
		214 =>	"00000100",	-- .....#..
		215 =>	"00000000",	-- ........

		-- char 0x1b='\x1b
		216 =>	"00000000",	-- ........
		217 =>	"00100000",	-- ..#.....
		218 =>	"01100000",	-- .##.....
		219 =>	"11111111",	-- ########
		220 =>	"11111111",	-- ########
		221 =>	"01100000",	-- .##.....
		222 =>	"00100000",	-- ..#.....
		223 =>	"00000000",	-- ........

		-- char 0x1c='\x1c
		224 =>	"00000000",	-- ........
		225 =>	"00000000",	-- ........
		226 =>	"11000000",	-- ##......
		227 =>	"11000000",	-- ##......
		228 =>	"11000000",	-- ##......
		229 =>	"11111110",	-- #######.
		230 =>	"00000000",	-- ........
		231 =>	"00000000",	-- ........

		-- char 0x1d='\x1d
		232 =>	"00000000",	-- ........
		233 =>	"00100100",	-- ..#..#..
		234 =>	"01100110",	-- .##..##.
		235 =>	"11111111",	-- ########
		236 =>	"11111111",	-- ########
		237 =>	"01100110",	-- .##..##.
		238 =>	"00100100",	-- ..#..#..
		239 =>	"00000000",	-- ........

		-- char 0x1e='\x1e
		240 =>	"00011000",	-- ...##...
		241 =>	"00011000",	-- ...##...
		242 =>	"00111100",	-- ..####..
		243 =>	"00111100",	-- ..####..
		244 =>	"01111110",	-- .######.
		245 =>	"01111110",	-- .######.
		246 =>	"11111111",	-- ########
		247 =>	"11111111",	-- ########

		-- char 0x1f='\x1f
		248 =>	"11111111",	-- ########
		249 =>	"11111111",	-- ########
		250 =>	"01111110",	-- .######.
		251 =>	"01111110",	-- .######.
		252 =>	"00111100",	-- ..####..
		253 =>	"00111100",	-- ..####..
		254 =>	"00011000",	-- ...##...
		255 =>	"00011000",	-- ...##...

		-- char 0x20=' '  
		256 =>	"00000000",	-- ........
		257 =>	"00000000",	-- ........
		258 =>	"00000000",	-- ........
		259 =>	"00000000",	-- ........
		260 =>	"00000000",	-- ........
		261 =>	"00000000",	-- ........
		262 =>	"00000000",	-- ........
		263 =>	"00000000",	-- ........

		-- char 0x21='!'  
		264 =>	"00110000",	-- ..##....
		265 =>	"01111000",	-- .####...
		266 =>	"01111000",	-- .####...
		267 =>	"00110000",	-- ..##....
		268 =>	"00110000",	-- ..##....
		269 =>	"00000000",	-- ........
		270 =>	"00110000",	-- ..##....
		271 =>	"00000000",	-- ........

		-- char 0x22='\'' 
		272 =>	"01101100",	-- .##.##..
		273 =>	"01101100",	-- .##.##..
		274 =>	"01101100",	-- .##.##..
		275 =>	"00000000",	-- ........
		276 =>	"00000000",	-- ........
		277 =>	"00000000",	-- ........
		278 =>	"00000000",	-- ........
		279 =>	"00000000",	-- ........

		-- char 0x23='#'  
		280 =>	"01101100",	-- .##.##..
		281 =>	"01101100",	-- .##.##..
		282 =>	"11111110",	-- #######.
		283 =>	"01101100",	-- .##.##..
		284 =>	"11111110",	-- #######.
		285 =>	"01101100",	-- .##.##..
		286 =>	"01101100",	-- .##.##..
		287 =>	"00000000",	-- ........

		-- char 0x24='$'  
		288 =>	"00110000",	-- ..##....
		289 =>	"01111100",	-- .#####..
		290 =>	"11000000",	-- ##......
		291 =>	"01111000",	-- .####...
		292 =>	"00001100",	-- ....##..
		293 =>	"11111000",	-- #####...
		294 =>	"00110000",	-- ..##....
		295 =>	"00000000",	-- ........

		-- char 0x25='%'  
		296 =>	"00000000",	-- ........
		297 =>	"11000110",	-- ##...##.
		298 =>	"11001100",	-- ##..##..
		299 =>	"00011000",	-- ...##...
		300 =>	"00110000",	-- ..##....
		301 =>	"01100110",	-- .##..##.
		302 =>	"11000110",	-- ##...##.
		303 =>	"00000000",	-- ........

		-- char 0x26='&'  
		304 =>	"00111000",	-- ..###...
		305 =>	"01101100",	-- .##.##..
		306 =>	"00111000",	-- ..###...
		307 =>	"01110110",	-- .###.##.
		308 =>	"11011100",	-- ##.###..
		309 =>	"11001100",	-- ##..##..
		310 =>	"01110110",	-- .###.##.
		311 =>	"00000000",	-- ........

		-- char 0x27='\"' 
		312 =>	"01100000",	-- .##.....
		313 =>	"01100000",	-- .##.....
		314 =>	"11000000",	-- ##......
		315 =>	"00000000",	-- ........
		316 =>	"00000000",	-- ........
		317 =>	"00000000",	-- ........
		318 =>	"00000000",	-- ........
		319 =>	"00000000",	-- ........

		-- char 0x28='('  
		320 =>	"00011000",	-- ...##...
		321 =>	"00110000",	-- ..##....
		322 =>	"01100000",	-- .##.....
		323 =>	"01100000",	-- .##.....
		324 =>	"01100000",	-- .##.....
		325 =>	"00110000",	-- ..##....
		326 =>	"00011000",	-- ...##...
		327 =>	"00000000",	-- ........

		-- char 0x29=')'  
		328 =>	"01100000",	-- .##.....
		329 =>	"00110000",	-- ..##....
		330 =>	"00011000",	-- ...##...
		331 =>	"00011000",	-- ...##...
		332 =>	"00011000",	-- ...##...
		333 =>	"00110000",	-- ..##....
		334 =>	"01100000",	-- .##.....
		335 =>	"00000000",	-- ........

		-- char 0x2a='*'  
		336 =>	"00000000",	-- ........
		337 =>	"01100110",	-- .##..##.
		338 =>	"00111100",	-- ..####..
		339 =>	"11111111",	-- ########
		340 =>	"00111100",	-- ..####..
		341 =>	"01100110",	-- .##..##.
		342 =>	"00000000",	-- ........
		343 =>	"00000000",	-- ........

		-- char 0x2b='+'  
		344 =>	"00000000",	-- ........
		345 =>	"00110000",	-- ..##....
		346 =>	"00110000",	-- ..##....
		347 =>	"11111100",	-- ######..
		348 =>	"00110000",	-- ..##....
		349 =>	"00110000",	-- ..##....
		350 =>	"00000000",	-- ........
		351 =>	"00000000",	-- ........

		-- char 0x2c=','  
		352 =>	"00000000",	-- ........
		353 =>	"00000000",	-- ........
		354 =>	"00000000",	-- ........
		355 =>	"00000000",	-- ........
		356 =>	"00000000",	-- ........
		357 =>	"01110000",	-- .###....
		358 =>	"00110000",	-- ..##....
		359 =>	"01100000",	-- .##.....

		-- char 0x2d='-'  
		360 =>	"00000000",	-- ........
		361 =>	"00000000",	-- ........
		362 =>	"00000000",	-- ........
		363 =>	"11111100",	-- ######..
		364 =>	"00000000",	-- ........
		365 =>	"00000000",	-- ........
		366 =>	"00000000",	-- ........
		367 =>	"00000000",	-- ........

		-- char 0x2e='.'  
		368 =>	"00000000",	-- ........
		369 =>	"00000000",	-- ........
		370 =>	"00000000",	-- ........
		371 =>	"00000000",	-- ........
		372 =>	"00000000",	-- ........
		373 =>	"00110000",	-- ..##....
		374 =>	"00110000",	-- ..##....
		375 =>	"00000000",	-- ........

		-- char 0x2f='/'  
		376 =>	"00000011",	-- ......##
		377 =>	"00000111",	-- .....###
		378 =>	"00001110",	-- ....###.
		379 =>	"00011100",	-- ...###..
		380 =>	"00111000",	-- ..###...
		381 =>	"01110000",	-- .###....
		382 =>	"11100000",	-- ###.....
		383 =>	"11000000",	-- ##......

		-- char 0x30='0'  
		384 =>	"01111000",	-- .####...
		385 =>	"11001100",	-- ##..##..
		386 =>	"11011100",	-- ##.###..
		387 =>	"11111100",	-- ######..
		388 =>	"11101100",	-- ###.##..
		389 =>	"11001100",	-- ##..##..
		390 =>	"01111000",	-- .####...
		391 =>	"00000000",	-- ........

		-- char 0x31='1'  
		392 =>	"00110000",	-- ..##....
		393 =>	"11110000",	-- ####....
		394 =>	"00110000",	-- ..##....
		395 =>	"00110000",	-- ..##....
		396 =>	"00110000",	-- ..##....
		397 =>	"00110000",	-- ..##....
		398 =>	"11111100",	-- ######..
		399 =>	"00000000",	-- ........

		-- char 0x32='2'  
		400 =>	"01111000",	-- .####...
		401 =>	"11001100",	-- ##..##..
		402 =>	"00001100",	-- ....##..
		403 =>	"00111000",	-- ..###...
		404 =>	"01100000",	-- .##.....
		405 =>	"11001100",	-- ##..##..
		406 =>	"11111100",	-- ######..
		407 =>	"00000000",	-- ........

		-- char 0x33='3'  
		408 =>	"01111000",	-- .####...
		409 =>	"11001100",	-- ##..##..
		410 =>	"00001100",	-- ....##..
		411 =>	"00111000",	-- ..###...
		412 =>	"00001100",	-- ....##..
		413 =>	"11001100",	-- ##..##..
		414 =>	"01111000",	-- .####...
		415 =>	"00000000",	-- ........

		-- char 0x34='4'  
		416 =>	"00011100",	-- ...###..
		417 =>	"00111100",	-- ..####..
		418 =>	"01101100",	-- .##.##..
		419 =>	"11001100",	-- ##..##..
		420 =>	"11111110",	-- #######.
		421 =>	"00001100",	-- ....##..
		422 =>	"00001100",	-- ....##..
		423 =>	"00000000",	-- ........

		-- char 0x35='5'  
		424 =>	"11111100",	-- ######..
		425 =>	"11000000",	-- ##......
		426 =>	"11111000",	-- #####...
		427 =>	"00001100",	-- ....##..
		428 =>	"00001100",	-- ....##..
		429 =>	"11001100",	-- ##..##..
		430 =>	"01111000",	-- .####...
		431 =>	"00000000",	-- ........

		-- char 0x36='6'  
		432 =>	"00111000",	-- ..###...
		433 =>	"01100000",	-- .##.....
		434 =>	"11000000",	-- ##......
		435 =>	"11111000",	-- #####...
		436 =>	"11001100",	-- ##..##..
		437 =>	"11001100",	-- ##..##..
		438 =>	"01111000",	-- .####...
		439 =>	"00000000",	-- ........

		-- char 0x37='7'  
		440 =>	"11111100",	-- ######..
		441 =>	"11001100",	-- ##..##..
		442 =>	"00001100",	-- ....##..
		443 =>	"00011000",	-- ...##...
		444 =>	"00110000",	-- ..##....
		445 =>	"01100000",	-- .##.....
		446 =>	"01100000",	-- .##.....
		447 =>	"00000000",	-- ........

		-- char 0x38='8'  
		448 =>	"01111000",	-- .####...
		449 =>	"11001100",	-- ##..##..
		450 =>	"11001100",	-- ##..##..
		451 =>	"01111000",	-- .####...
		452 =>	"11001100",	-- ##..##..
		453 =>	"11001100",	-- ##..##..
		454 =>	"01111000",	-- .####...
		455 =>	"00000000",	-- ........

		-- char 0x39='9'  
		456 =>	"01111000",	-- .####...
		457 =>	"11001100",	-- ##..##..
		458 =>	"11001100",	-- ##..##..
		459 =>	"01111100",	-- .#####..
		460 =>	"00001100",	-- ....##..
		461 =>	"00011000",	-- ...##...
		462 =>	"01110000",	-- .###....
		463 =>	"00000000",	-- ........

		-- char 0x3a=':'  
		464 =>	"00000000",	-- ........
		465 =>	"00000000",	-- ........
		466 =>	"00110000",	-- ..##....
		467 =>	"00110000",	-- ..##....
		468 =>	"00000000",	-- ........
		469 =>	"00110000",	-- ..##....
		470 =>	"00110000",	-- ..##....
		471 =>	"00000000",	-- ........

		-- char 0x3b=';'  
		472 =>	"00000000",	-- ........
		473 =>	"00000000",	-- ........
		474 =>	"00110000",	-- ..##....
		475 =>	"00110000",	-- ..##....
		476 =>	"00000000",	-- ........
		477 =>	"01110000",	-- .###....
		478 =>	"00110000",	-- ..##....
		479 =>	"01100000",	-- .##.....

		-- char 0x3c='<'  
		480 =>	"00011000",	-- ...##...
		481 =>	"00110000",	-- ..##....
		482 =>	"01100000",	-- .##.....
		483 =>	"11000000",	-- ##......
		484 =>	"01100000",	-- .##.....
		485 =>	"00110000",	-- ..##....
		486 =>	"00011000",	-- ...##...
		487 =>	"00000000",	-- ........

		-- char 0x3d='='  
		488 =>	"00000000",	-- ........
		489 =>	"00000000",	-- ........
		490 =>	"11111100",	-- ######..
		491 =>	"00000000",	-- ........
		492 =>	"11111100",	-- ######..
		493 =>	"00000000",	-- ........
		494 =>	"00000000",	-- ........
		495 =>	"00000000",	-- ........

		-- char 0x3e='>'  
		496 =>	"01100000",	-- .##.....
		497 =>	"00110000",	-- ..##....
		498 =>	"00011000",	-- ...##...
		499 =>	"00001100",	-- ....##..
		500 =>	"00011000",	-- ...##...
		501 =>	"00110000",	-- ..##....
		502 =>	"01100000",	-- .##.....
		503 =>	"00000000",	-- ........

		-- char 0x3f='?'  
		504 =>	"01111000",	-- .####...
		505 =>	"11001100",	-- ##..##..
		506 =>	"00001100",	-- ....##..
		507 =>	"00011000",	-- ...##...
		508 =>	"00110000",	-- ..##....
		509 =>	"00000000",	-- ........
		510 =>	"00110000",	-- ..##....
		511 =>	"00000000",	-- ........

		-- char 0x40='@'  
		512 =>	"01111100",	-- .#####..
		513 =>	"11000110",	-- ##...##.
		514 =>	"11011110",	-- ##.####.
		515 =>	"11011110",	-- ##.####.
		516 =>	"11011110",	-- ##.####.
		517 =>	"11000000",	-- ##......
		518 =>	"01111000",	-- .####...
		519 =>	"00000000",	-- ........

		-- char 0x41='A'  
		520 =>	"00110000",	-- ..##....
		521 =>	"01111000",	-- .####...
		522 =>	"11001100",	-- ##..##..
		523 =>	"11001100",	-- ##..##..
		524 =>	"11111100",	-- ######..
		525 =>	"11001100",	-- ##..##..
		526 =>	"11001100",	-- ##..##..
		527 =>	"00000000",	-- ........

		-- char 0x42='B'  
		528 =>	"11111100",	-- ######..
		529 =>	"01100110",	-- .##..##.
		530 =>	"01100110",	-- .##..##.
		531 =>	"01111100",	-- .#####..
		532 =>	"01100110",	-- .##..##.
		533 =>	"01100110",	-- .##..##.
		534 =>	"11111100",	-- ######..
		535 =>	"00000000",	-- ........

		-- char 0x43='C'  
		536 =>	"00111100",	-- ..####..
		537 =>	"01100110",	-- .##..##.
		538 =>	"11000000",	-- ##......
		539 =>	"11000000",	-- ##......
		540 =>	"11000000",	-- ##......
		541 =>	"01100110",	-- .##..##.
		542 =>	"00111100",	-- ..####..
		543 =>	"00000000",	-- ........

		-- char 0x44='D'  
		544 =>	"11111100",	-- ######..
		545 =>	"01101100",	-- .##.##..
		546 =>	"01100110",	-- .##..##.
		547 =>	"01100110",	-- .##..##.
		548 =>	"01100110",	-- .##..##.
		549 =>	"01101100",	-- .##.##..
		550 =>	"11111100",	-- ######..
		551 =>	"00000000",	-- ........

		-- char 0x45='E'  
		552 =>	"11111110",	-- #######.
		553 =>	"01100010",	-- .##...#.
		554 =>	"01101000",	-- .##.#...
		555 =>	"01111000",	-- .####...
		556 =>	"01101000",	-- .##.#...
		557 =>	"01100010",	-- .##...#.
		558 =>	"11111110",	-- #######.
		559 =>	"00000000",	-- ........

		-- char 0x46='F'  
		560 =>	"11111110",	-- #######.
		561 =>	"01100010",	-- .##...#.
		562 =>	"01101000",	-- .##.#...
		563 =>	"01111000",	-- .####...
		564 =>	"01101000",	-- .##.#...
		565 =>	"01100000",	-- .##.....
		566 =>	"11110000",	-- ####....
		567 =>	"00000000",	-- ........

		-- char 0x47='G'  
		568 =>	"00111100",	-- ..####..
		569 =>	"01100110",	-- .##..##.
		570 =>	"11000000",	-- ##......
		571 =>	"11000000",	-- ##......
		572 =>	"11001110",	-- ##..###.
		573 =>	"01100110",	-- .##..##.
		574 =>	"00111110",	-- ..#####.
		575 =>	"00000000",	-- ........

		-- char 0x48='H'  
		576 =>	"11001100",	-- ##..##..
		577 =>	"11001100",	-- ##..##..
		578 =>	"11001100",	-- ##..##..
		579 =>	"11111100",	-- ######..
		580 =>	"11001100",	-- ##..##..
		581 =>	"11001100",	-- ##..##..
		582 =>	"11001100",	-- ##..##..
		583 =>	"00000000",	-- ........

		-- char 0x49='I'  
		584 =>	"01111000",	-- .####...
		585 =>	"00110000",	-- ..##....
		586 =>	"00110000",	-- ..##....
		587 =>	"00110000",	-- ..##....
		588 =>	"00110000",	-- ..##....
		589 =>	"00110000",	-- ..##....
		590 =>	"01111000",	-- .####...
		591 =>	"00000000",	-- ........

		-- char 0x4a='J'  
		592 =>	"00011110",	-- ...####.
		593 =>	"00001100",	-- ....##..
		594 =>	"00001100",	-- ....##..
		595 =>	"00001100",	-- ....##..
		596 =>	"11001100",	-- ##..##..
		597 =>	"11001100",	-- ##..##..
		598 =>	"01111000",	-- .####...
		599 =>	"00000000",	-- ........

		-- char 0x4b='K'  
		600 =>	"11100110",	-- ###..##.
		601 =>	"01100110",	-- .##..##.
		602 =>	"01101100",	-- .##.##..
		603 =>	"01111000",	-- .####...
		604 =>	"01101100",	-- .##.##..
		605 =>	"01100110",	-- .##..##.
		606 =>	"11100110",	-- ###..##.
		607 =>	"00000000",	-- ........

		-- char 0x4c='L'  
		608 =>	"11110000",	-- ####....
		609 =>	"01100000",	-- .##.....
		610 =>	"01100000",	-- .##.....
		611 =>	"01100000",	-- .##.....
		612 =>	"01100010",	-- .##...#.
		613 =>	"01100110",	-- .##..##.
		614 =>	"11111110",	-- #######.
		615 =>	"00000000",	-- ........

		-- char 0x4d='M'  
		616 =>	"11000110",	-- ##...##.
		617 =>	"11101110",	-- ###.###.
		618 =>	"11111110",	-- #######.
		619 =>	"11010110",	-- ##.#.##.
		620 =>	"11000110",	-- ##...##.
		621 =>	"11000110",	-- ##...##.
		622 =>	"11000110",	-- ##...##.
		623 =>	"00000000",	-- ........

		-- char 0x4e='N'  
		624 =>	"11000110",	-- ##...##.
		625 =>	"11100110",	-- ###..##.
		626 =>	"11110110",	-- ####.##.
		627 =>	"11011110",	-- ##.####.
		628 =>	"11001110",	-- ##..###.
		629 =>	"11000110",	-- ##...##.
		630 =>	"11000110",	-- ##...##.
		631 =>	"00000000",	-- ........

		-- char 0x4f='O'  
		632 =>	"00111000",	-- ..###...
		633 =>	"01101100",	-- .##.##..
		634 =>	"11000110",	-- ##...##.
		635 =>	"11000110",	-- ##...##.
		636 =>	"11000110",	-- ##...##.
		637 =>	"01101100",	-- .##.##..
		638 =>	"00111000",	-- ..###...
		639 =>	"00000000",	-- ........

		-- char 0x50='P'  
		640 =>	"11111100",	-- ######..
		641 =>	"01100110",	-- .##..##.
		642 =>	"01100110",	-- .##..##.
		643 =>	"01111100",	-- .#####..
		644 =>	"01100000",	-- .##.....
		645 =>	"01100000",	-- .##.....
		646 =>	"11110000",	-- ####....
		647 =>	"00000000",	-- ........

		-- char 0x51='Q'  
		648 =>	"01111000",	-- .####...
		649 =>	"11001100",	-- ##..##..
		650 =>	"11001100",	-- ##..##..
		651 =>	"11001100",	-- ##..##..
		652 =>	"11011100",	-- ##.###..
		653 =>	"01111000",	-- .####...
		654 =>	"00011100",	-- ...###..
		655 =>	"00000000",	-- ........

		-- char 0x52='R'  
		656 =>	"11111100",	-- ######..
		657 =>	"01100110",	-- .##..##.
		658 =>	"01100110",	-- .##..##.
		659 =>	"01111100",	-- .#####..
		660 =>	"01111000",	-- .####...
		661 =>	"01101100",	-- .##.##..
		662 =>	"11100110",	-- ###..##.
		663 =>	"00000000",	-- ........

		-- char 0x53='S'  
		664 =>	"01111000",	-- .####...
		665 =>	"11001100",	-- ##..##..
		666 =>	"11100000",	-- ###.....
		667 =>	"00111000",	-- ..###...
		668 =>	"00011100",	-- ...###..
		669 =>	"11001100",	-- ##..##..
		670 =>	"01111000",	-- .####...
		671 =>	"00000000",	-- ........

		-- char 0x54='T'  
		672 =>	"11111100",	-- ######..
		673 =>	"10110100",	-- #.##.#..
		674 =>	"00110000",	-- ..##....
		675 =>	"00110000",	-- ..##....
		676 =>	"00110000",	-- ..##....
		677 =>	"00110000",	-- ..##....
		678 =>	"01111000",	-- .####...
		679 =>	"00000000",	-- ........

		-- char 0x55='U'  
		680 =>	"11001100",	-- ##..##..
		681 =>	"11001100",	-- ##..##..
		682 =>	"11001100",	-- ##..##..
		683 =>	"11001100",	-- ##..##..
		684 =>	"11001100",	-- ##..##..
		685 =>	"11001100",	-- ##..##..
		686 =>	"11111100",	-- ######..
		687 =>	"00000000",	-- ........

		-- char 0x56='V'  
		688 =>	"11001100",	-- ##..##..
		689 =>	"11001100",	-- ##..##..
		690 =>	"11001100",	-- ##..##..
		691 =>	"11001100",	-- ##..##..
		692 =>	"11001100",	-- ##..##..
		693 =>	"01111000",	-- .####...
		694 =>	"00110000",	-- ..##....
		695 =>	"00000000",	-- ........

		-- char 0x57='W'  
		696 =>	"11000110",	-- ##...##.
		697 =>	"11000110",	-- ##...##.
		698 =>	"11000110",	-- ##...##.
		699 =>	"11010110",	-- ##.#.##.
		700 =>	"11111110",	-- #######.
		701 =>	"11101110",	-- ###.###.
		702 =>	"11000110",	-- ##...##.
		703 =>	"00000000",	-- ........

		-- char 0x58='X'  
		704 =>	"11000110",	-- ##...##.
		705 =>	"11000110",	-- ##...##.
		706 =>	"01101100",	-- .##.##..
		707 =>	"00111000",	-- ..###...
		708 =>	"01101100",	-- .##.##..
		709 =>	"11000110",	-- ##...##.
		710 =>	"11000110",	-- ##...##.
		711 =>	"00000000",	-- ........

		-- char 0x59='Y'  
		712 =>	"11001100",	-- ##..##..
		713 =>	"11001100",	-- ##..##..
		714 =>	"11001100",	-- ##..##..
		715 =>	"01111000",	-- .####...
		716 =>	"00110000",	-- ..##....
		717 =>	"00110000",	-- ..##....
		718 =>	"01111000",	-- .####...
		719 =>	"00000000",	-- ........

		-- char 0x5a='Z'  
		720 =>	"11111110",	-- #######.
		721 =>	"11001100",	-- ##..##..
		722 =>	"10011000",	-- #..##...
		723 =>	"00110000",	-- ..##....
		724 =>	"01100010",	-- .##...#.
		725 =>	"11000110",	-- ##...##.
		726 =>	"11111110",	-- #######.
		727 =>	"00000000",	-- ........

		-- char 0x5b='['  
		728 =>	"01111000",	-- .####...
		729 =>	"01100000",	-- .##.....
		730 =>	"01100000",	-- .##.....
		731 =>	"01100000",	-- .##.....
		732 =>	"01100000",	-- .##.....
		733 =>	"01100000",	-- .##.....
		734 =>	"01111000",	-- .####...
		735 =>	"00000000",	-- ........

		-- char 0x5c='\\' 
		736 =>	"11000000",	-- ##......
		737 =>	"11100000",	-- ###.....
		738 =>	"01110000",	-- .###....
		739 =>	"00111000",	-- ..###...
		740 =>	"00011100",	-- ...###..
		741 =>	"00001110",	-- ....###.
		742 =>	"00000111",	-- .....###
		743 =>	"00000011",	-- ......##

		-- char 0x5d=']'  
		744 =>	"01111000",	-- .####...
		745 =>	"00011000",	-- ...##...
		746 =>	"00011000",	-- ...##...
		747 =>	"00011000",	-- ...##...
		748 =>	"00011000",	-- ...##...
		749 =>	"00011000",	-- ...##...
		750 =>	"01111000",	-- .####...
		751 =>	"00000000",	-- ........

		-- char 0x5e='^'  
		752 =>	"00010000",	-- ...#....
		753 =>	"00111000",	-- ..###...
		754 =>	"01101100",	-- .##.##..
		755 =>	"11000110",	-- ##...##.
		756 =>	"00000000",	-- ........
		757 =>	"00000000",	-- ........
		758 =>	"00000000",	-- ........
		759 =>	"00000000",	-- ........

		-- char 0x5f='_'  
		760 =>	"00000000",	-- ........
		761 =>	"00000000",	-- ........
		762 =>	"00000000",	-- ........
		763 =>	"00000000",	-- ........
		764 =>	"00000000",	-- ........
		765 =>	"00000000",	-- ........
		766 =>	"00000000",	-- ........
		767 =>	"11111111",	-- ########

		-- char 0x60='`'  
		768 =>	"00110000",	-- ..##....
		769 =>	"00110000",	-- ..##....
		770 =>	"00011000",	-- ...##...
		771 =>	"00000000",	-- ........
		772 =>	"00000000",	-- ........
		773 =>	"00000000",	-- ........
		774 =>	"00000000",	-- ........
		775 =>	"00000000",	-- ........

		-- char 0x61='a'  
		776 =>	"00000000",	-- ........
		777 =>	"00000000",	-- ........
		778 =>	"01111000",	-- .####...
		779 =>	"00001100",	-- ....##..
		780 =>	"01111100",	-- .#####..
		781 =>	"11001100",	-- ##..##..
		782 =>	"01110110",	-- .###.##.
		783 =>	"00000000",	-- ........

		-- char 0x62='b'  
		784 =>	"11100000",	-- ###.....
		785 =>	"01100000",	-- .##.....
		786 =>	"01111100",	-- .#####..
		787 =>	"01100110",	-- .##..##.
		788 =>	"01100110",	-- .##..##.
		789 =>	"01100110",	-- .##..##.
		790 =>	"10111100",	-- #.####..
		791 =>	"00000000",	-- ........

		-- char 0x63='c'  
		792 =>	"00000000",	-- ........
		793 =>	"00000000",	-- ........
		794 =>	"01111000",	-- .####...
		795 =>	"11001100",	-- ##..##..
		796 =>	"11000000",	-- ##......
		797 =>	"11001100",	-- ##..##..
		798 =>	"01111000",	-- .####...
		799 =>	"00000000",	-- ........

		-- char 0x64='d'  
		800 =>	"00011100",	-- ...###..
		801 =>	"00001100",	-- ....##..
		802 =>	"00001100",	-- ....##..
		803 =>	"01111100",	-- .#####..
		804 =>	"11001100",	-- ##..##..
		805 =>	"11001100",	-- ##..##..
		806 =>	"01110110",	-- .###.##.
		807 =>	"00000000",	-- ........

		-- char 0x65='e'  
		808 =>	"00000000",	-- ........
		809 =>	"00000000",	-- ........
		810 =>	"01111000",	-- .####...
		811 =>	"11001100",	-- ##..##..
		812 =>	"11111100",	-- ######..
		813 =>	"11000000",	-- ##......
		814 =>	"01111000",	-- .####...
		815 =>	"00000000",	-- ........

		-- char 0x66='f'  
		816 =>	"00111000",	-- ..###...
		817 =>	"01101100",	-- .##.##..
		818 =>	"01100000",	-- .##.....
		819 =>	"11110000",	-- ####....
		820 =>	"01100000",	-- .##.....
		821 =>	"01100000",	-- .##.....
		822 =>	"11110000",	-- ####....
		823 =>	"00000000",	-- ........

		-- char 0x67='g'  
		824 =>	"00000000",	-- ........
		825 =>	"00000000",	-- ........
		826 =>	"01110110",	-- .###.##.
		827 =>	"11001100",	-- ##..##..
		828 =>	"11001100",	-- ##..##..
		829 =>	"01111100",	-- .#####..
		830 =>	"00001100",	-- ....##..
		831 =>	"11111000",	-- #####...

		-- char 0x68='h'  
		832 =>	"11100000",	-- ###.....
		833 =>	"01100000",	-- .##.....
		834 =>	"01101100",	-- .##.##..
		835 =>	"01110110",	-- .###.##.
		836 =>	"01100110",	-- .##..##.
		837 =>	"01100110",	-- .##..##.
		838 =>	"11100110",	-- ###..##.
		839 =>	"00000000",	-- ........

		-- char 0x69='i'  
		840 =>	"00110000",	-- ..##....
		841 =>	"00000000",	-- ........
		842 =>	"01110000",	-- .###....
		843 =>	"00110000",	-- ..##....
		844 =>	"00110000",	-- ..##....
		845 =>	"00110000",	-- ..##....
		846 =>	"01111000",	-- .####...
		847 =>	"00000000",	-- ........

		-- char 0x6a='j'  
		848 =>	"00011000",	-- ...##...
		849 =>	"00000000",	-- ........
		850 =>	"01111000",	-- .####...
		851 =>	"00011000",	-- ...##...
		852 =>	"00011000",	-- ...##...
		853 =>	"00011000",	-- ...##...
		854 =>	"11011000",	-- ##.##...
		855 =>	"01110000",	-- .###....

		-- char 0x6b='k'  
		856 =>	"11100000",	-- ###.....
		857 =>	"01100000",	-- .##.....
		858 =>	"01100110",	-- .##..##.
		859 =>	"01101100",	-- .##.##..
		860 =>	"01111000",	-- .####...
		861 =>	"01101100",	-- .##.##..
		862 =>	"11100110",	-- ###..##.
		863 =>	"00000000",	-- ........

		-- char 0x6c='l'  
		864 =>	"01110000",	-- .###....
		865 =>	"00110000",	-- ..##....
		866 =>	"00110000",	-- ..##....
		867 =>	"00110000",	-- ..##....
		868 =>	"00110000",	-- ..##....
		869 =>	"00110000",	-- ..##....
		870 =>	"01111000",	-- .####...
		871 =>	"00000000",	-- ........

		-- char 0x6d='m'  
		872 =>	"00000000",	-- ........
		873 =>	"00000000",	-- ........
		874 =>	"11101100",	-- ###.##..
		875 =>	"11111110",	-- #######.
		876 =>	"11010110",	-- ##.#.##.
		877 =>	"11000110",	-- ##...##.
		878 =>	"11000110",	-- ##...##.
		879 =>	"00000000",	-- ........

		-- char 0x6e='n'  
		880 =>	"00000000",	-- ........
		881 =>	"00000000",	-- ........
		882 =>	"11111000",	-- #####...
		883 =>	"11001100",	-- ##..##..
		884 =>	"11001100",	-- ##..##..
		885 =>	"11001100",	-- ##..##..
		886 =>	"11001100",	-- ##..##..
		887 =>	"00000000",	-- ........

		-- char 0x6f='o'  
		888 =>	"00000000",	-- ........
		889 =>	"00000000",	-- ........
		890 =>	"01111000",	-- .####...
		891 =>	"11001100",	-- ##..##..
		892 =>	"11001100",	-- ##..##..
		893 =>	"11001100",	-- ##..##..
		894 =>	"01111000",	-- .####...
		895 =>	"00000000",	-- ........

		-- char 0x70='p'  
		896 =>	"00000000",	-- ........
		897 =>	"00000000",	-- ........
		898 =>	"11011100",	-- ##.###..
		899 =>	"01100110",	-- .##..##.
		900 =>	"01100110",	-- .##..##.
		901 =>	"01111100",	-- .#####..
		902 =>	"01100000",	-- .##.....
		903 =>	"11110000",	-- ####....

		-- char 0x71='q'  
		904 =>	"00000000",	-- ........
		905 =>	"00000000",	-- ........
		906 =>	"01110110",	-- .###.##.
		907 =>	"11001100",	-- ##..##..
		908 =>	"11001100",	-- ##..##..
		909 =>	"01111100",	-- .#####..
		910 =>	"00001100",	-- ....##..
		911 =>	"00011110",	-- ...####.

		-- char 0x72='r'  
		912 =>	"00000000",	-- ........
		913 =>	"00000000",	-- ........
		914 =>	"11011000",	-- ##.##...
		915 =>	"01101100",	-- .##.##..
		916 =>	"01101100",	-- .##.##..
		917 =>	"01100000",	-- .##.....
		918 =>	"11110000",	-- ####....
		919 =>	"00000000",	-- ........

		-- char 0x73='s'  
		920 =>	"00000000",	-- ........
		921 =>	"00000000",	-- ........
		922 =>	"01111100",	-- .#####..
		923 =>	"11000000",	-- ##......
		924 =>	"01111000",	-- .####...
		925 =>	"00001100",	-- ....##..
		926 =>	"11111000",	-- #####...
		927 =>	"00000000",	-- ........

		-- char 0x74='t'  
		928 =>	"00010000",	-- ...#....
		929 =>	"00110000",	-- ..##....
		930 =>	"01111100",	-- .#####..
		931 =>	"00110000",	-- ..##....
		932 =>	"00110000",	-- ..##....
		933 =>	"00110100",	-- ..##.#..
		934 =>	"00011000",	-- ...##...
		935 =>	"00000000",	-- ........

		-- char 0x75='u'  
		936 =>	"00000000",	-- ........
		937 =>	"00000000",	-- ........
		938 =>	"11001100",	-- ##..##..
		939 =>	"11001100",	-- ##..##..
		940 =>	"11001100",	-- ##..##..
		941 =>	"11001100",	-- ##..##..
		942 =>	"01110110",	-- .###.##.
		943 =>	"00000000",	-- ........

		-- char 0x76='v'  
		944 =>	"00000000",	-- ........
		945 =>	"00000000",	-- ........
		946 =>	"11001100",	-- ##..##..
		947 =>	"11001100",	-- ##..##..
		948 =>	"11001100",	-- ##..##..
		949 =>	"01111000",	-- .####...
		950 =>	"00110000",	-- ..##....
		951 =>	"00000000",	-- ........

		-- char 0x77='w'  
		952 =>	"00000000",	-- ........
		953 =>	"00000000",	-- ........
		954 =>	"11000110",	-- ##...##.
		955 =>	"11000110",	-- ##...##.
		956 =>	"11010110",	-- ##.#.##.
		957 =>	"11111110",	-- #######.
		958 =>	"01101100",	-- .##.##..
		959 =>	"00000000",	-- ........

		-- char 0x78='x'  
		960 =>	"00000000",	-- ........
		961 =>	"00000000",	-- ........
		962 =>	"11000110",	-- ##...##.
		963 =>	"01101100",	-- .##.##..
		964 =>	"00111000",	-- ..###...
		965 =>	"01101100",	-- .##.##..
		966 =>	"11000110",	-- ##...##.
		967 =>	"00000000",	-- ........

		-- char 0x79='y'  
		968 =>	"00000000",	-- ........
		969 =>	"00000000",	-- ........
		970 =>	"11001100",	-- ##..##..
		971 =>	"11001100",	-- ##..##..
		972 =>	"11001100",	-- ##..##..
		973 =>	"01111100",	-- .#####..
		974 =>	"00001100",	-- ....##..
		975 =>	"11111000",	-- #####...

		-- char 0x7a='z'  
		976 =>	"00000000",	-- ........
		977 =>	"00000000",	-- ........
		978 =>	"11111100",	-- ######..
		979 =>	"10011000",	-- #..##...
		980 =>	"00110000",	-- ..##....
		981 =>	"01100100",	-- .##..#..
		982 =>	"11111100",	-- ######..
		983 =>	"00000000",	-- ........

		-- char 0x7b='{'  
		984 =>	"00011100",	-- ...###..
		985 =>	"00110000",	-- ..##....
		986 =>	"00110000",	-- ..##....
		987 =>	"11100000",	-- ###.....
		988 =>	"00110000",	-- ..##....
		989 =>	"00110000",	-- ..##....
		990 =>	"00011100",	-- ...###..
		991 =>	"00000000",	-- ........

		-- char 0x7c='|'  
		992 =>	"00011000",	-- ...##...
		993 =>	"00011000",	-- ...##...
		994 =>	"00011000",	-- ...##...
		995 =>	"00000000",	-- ........
		996 =>	"00011000",	-- ...##...
		997 =>	"00011000",	-- ...##...
		998 =>	"00011000",	-- ...##...
		999 =>	"00000000",	-- ........

		-- char 0x7d='}'  
		1000 =>	"11100000",	-- ###.....
		1001 =>	"00110000",	-- ..##....
		1002 =>	"00110000",	-- ..##....
		1003 =>	"00011100",	-- ...###..
		1004 =>	"00110000",	-- ..##....
		1005 =>	"00110000",	-- ..##....
		1006 =>	"11100000",	-- ###.....
		1007 =>	"00000000",	-- ........

		-- char 0x7e='~'  
		1008 =>	"01110110",	-- .###.##.
		1009 =>	"11011100",	-- ##.###..
		1010 =>	"00000000",	-- ........
		1011 =>	"00000000",	-- ........
		1012 =>	"00000000",	-- ........
		1013 =>	"00000000",	-- ........
		1014 =>	"00000000",	-- ........
		1015 =>	"00000000",	-- ........

		-- char 0x7f='\x7f
		1016 =>	"00011000",	-- ...##...
		1017 =>	"00111100",	-- ..####..
		1018 =>	"01100110",	-- .##..##.
		1019 =>	"11000011",	-- ##....##
		1020 =>	"11000011",	-- ##....##
		1021 =>	"11000011",	-- ##....##
		1022 =>	"11000011",	-- ##....##
		1023 =>	"11111111",	-- ########

		-- char 0x80='\x80
		1024 =>	"01111000",	-- .####...
		1025 =>	"11001100",	-- ##..##..
		1026 =>	"11000000",	-- ##......
		1027 =>	"11000000",	-- ##......
		1028 =>	"11001100",	-- ##..##..
		1029 =>	"01111000",	-- .####...
		1030 =>	"00110000",	-- ..##....
		1031 =>	"01100000",	-- .##.....

		-- char 0x81='\x81
		1032 =>	"00000000",	-- ........
		1033 =>	"11001100",	-- ##..##..
		1034 =>	"00000000",	-- ........
		1035 =>	"11001100",	-- ##..##..
		1036 =>	"11001100",	-- ##..##..
		1037 =>	"11001100",	-- ##..##..
		1038 =>	"01111110",	-- .######.
		1039 =>	"00000000",	-- ........

		-- char 0x82='\x82
		1040 =>	"00011000",	-- ...##...
		1041 =>	"00110000",	-- ..##....
		1042 =>	"01111000",	-- .####...
		1043 =>	"11001100",	-- ##..##..
		1044 =>	"11111100",	-- ######..
		1045 =>	"11000000",	-- ##......
		1046 =>	"01111000",	-- .####...
		1047 =>	"00000000",	-- ........

		-- char 0x83='\x83
		1048 =>	"01111110",	-- .######.
		1049 =>	"11000011",	-- ##....##
		1050 =>	"00111100",	-- ..####..
		1051 =>	"00000110",	-- .....##.
		1052 =>	"00111110",	-- ..#####.
		1053 =>	"01100110",	-- .##..##.
		1054 =>	"00111111",	-- ..######
		1055 =>	"00000000",	-- ........

		-- char 0x84='\x84
		1056 =>	"11001100",	-- ##..##..
		1057 =>	"00000000",	-- ........
		1058 =>	"01111000",	-- .####...
		1059 =>	"00001100",	-- ....##..
		1060 =>	"01111100",	-- .#####..
		1061 =>	"11001100",	-- ##..##..
		1062 =>	"01111110",	-- .######.
		1063 =>	"00000000",	-- ........

		-- char 0x85='\x85
		1064 =>	"01100000",	-- .##.....
		1065 =>	"00110000",	-- ..##....
		1066 =>	"01111000",	-- .####...
		1067 =>	"00001100",	-- ....##..
		1068 =>	"01111100",	-- .#####..
		1069 =>	"11001100",	-- ##..##..
		1070 =>	"01111110",	-- .######.
		1071 =>	"00000000",	-- ........

		-- char 0x86='\x86
		1072 =>	"00111100",	-- ..####..
		1073 =>	"01100110",	-- .##..##.
		1074 =>	"00111100",	-- ..####..
		1075 =>	"00000110",	-- .....##.
		1076 =>	"00111110",	-- ..#####.
		1077 =>	"01100110",	-- .##..##.
		1078 =>	"00111111",	-- ..######
		1079 =>	"00000000",	-- ........

		-- char 0x87='\x87
		1080 =>	"00000000",	-- ........
		1081 =>	"01111000",	-- .####...
		1082 =>	"11001100",	-- ##..##..
		1083 =>	"11000000",	-- ##......
		1084 =>	"11001100",	-- ##..##..
		1085 =>	"01111000",	-- .####...
		1086 =>	"00110000",	-- ..##....
		1087 =>	"01100000",	-- .##.....

		-- char 0x88='\x88
		1088 =>	"01111110",	-- .######.
		1089 =>	"11000011",	-- ##....##
		1090 =>	"00111100",	-- ..####..
		1091 =>	"01100110",	-- .##..##.
		1092 =>	"01111110",	-- .######.
		1093 =>	"01100000",	-- .##.....
		1094 =>	"00111100",	-- ..####..
		1095 =>	"00000000",	-- ........

		-- char 0x89='\x89
		1096 =>	"11001100",	-- ##..##..
		1097 =>	"00000000",	-- ........
		1098 =>	"01111000",	-- .####...
		1099 =>	"11001100",	-- ##..##..
		1100 =>	"11111100",	-- ######..
		1101 =>	"11000000",	-- ##......
		1102 =>	"01111000",	-- .####...
		1103 =>	"00000000",	-- ........

		-- char 0x8a='\x8a
		1104 =>	"01100000",	-- .##.....
		1105 =>	"00110000",	-- ..##....
		1106 =>	"01111000",	-- .####...
		1107 =>	"11001100",	-- ##..##..
		1108 =>	"11111100",	-- ######..
		1109 =>	"11000000",	-- ##......
		1110 =>	"01111000",	-- .####...
		1111 =>	"00000000",	-- ........

		-- char 0x8b='\x8b
		1112 =>	"11001100",	-- ##..##..
		1113 =>	"00000000",	-- ........
		1114 =>	"01110000",	-- .###....
		1115 =>	"00110000",	-- ..##....
		1116 =>	"00110000",	-- ..##....
		1117 =>	"00110000",	-- ..##....
		1118 =>	"01111000",	-- .####...
		1119 =>	"00000000",	-- ........

		-- char 0x8c='\x8c
		1120 =>	"01111100",	-- .#####..
		1121 =>	"11000110",	-- ##...##.
		1122 =>	"00111000",	-- ..###...
		1123 =>	"00011000",	-- ...##...
		1124 =>	"00011000",	-- ...##...
		1125 =>	"00011000",	-- ...##...
		1126 =>	"00111100",	-- ..####..
		1127 =>	"00000000",	-- ........

		-- char 0x8d='\x8d
		1128 =>	"01100000",	-- .##.....
		1129 =>	"00110000",	-- ..##....
		1130 =>	"01110000",	-- .###....
		1131 =>	"00110000",	-- ..##....
		1132 =>	"00110000",	-- ..##....
		1133 =>	"00110000",	-- ..##....
		1134 =>	"01111000",	-- .####...
		1135 =>	"00000000",	-- ........

		-- char 0x8e='\x8e
		1136 =>	"11001100",	-- ##..##..
		1137 =>	"00110000",	-- ..##....
		1138 =>	"01111000",	-- .####...
		1139 =>	"11001100",	-- ##..##..
		1140 =>	"11001100",	-- ##..##..
		1141 =>	"11111100",	-- ######..
		1142 =>	"11001100",	-- ##..##..
		1143 =>	"00000000",	-- ........

		-- char 0x8f='\x8f
		1144 =>	"00110000",	-- ..##....
		1145 =>	"01001000",	-- .#..#...
		1146 =>	"00110000",	-- ..##....
		1147 =>	"01111000",	-- .####...
		1148 =>	"11001100",	-- ##..##..
		1149 =>	"11111100",	-- ######..
		1150 =>	"11001100",	-- ##..##..
		1151 =>	"00000000",	-- ........

		-- char 0x90='\x90
		1152 =>	"00011000",	-- ...##...
		1153 =>	"00110000",	-- ..##....
		1154 =>	"11111100",	-- ######..
		1155 =>	"01100000",	-- .##.....
		1156 =>	"01111000",	-- .####...
		1157 =>	"01100000",	-- .##.....
		1158 =>	"11111100",	-- ######..
		1159 =>	"00000000",	-- ........

		-- char 0x91='\x91
		1160 =>	"00000000",	-- ........
		1161 =>	"00000000",	-- ........
		1162 =>	"01111111",	-- .#######
		1163 =>	"00001100",	-- ....##..
		1164 =>	"01111111",	-- .#######
		1165 =>	"11001100",	-- ##..##..
		1166 =>	"01111111",	-- .#######
		1167 =>	"00000000",	-- ........

		-- char 0x92='\x92
		1168 =>	"00111110",	-- ..#####.
		1169 =>	"01101100",	-- .##.##..
		1170 =>	"11001100",	-- ##..##..
		1171 =>	"11111110",	-- #######.
		1172 =>	"11001100",	-- ##..##..
		1173 =>	"11001100",	-- ##..##..
		1174 =>	"11001110",	-- ##..###.
		1175 =>	"00000000",	-- ........

		-- char 0x93='\x93
		1176 =>	"01111000",	-- .####...
		1177 =>	"11001100",	-- ##..##..
		1178 =>	"00000000",	-- ........
		1179 =>	"01111000",	-- .####...
		1180 =>	"11001100",	-- ##..##..
		1181 =>	"11001100",	-- ##..##..
		1182 =>	"01111000",	-- .####...
		1183 =>	"00000000",	-- ........

		-- char 0x94='\x94
		1184 =>	"00000000",	-- ........
		1185 =>	"11001100",	-- ##..##..
		1186 =>	"00000000",	-- ........
		1187 =>	"01111000",	-- .####...
		1188 =>	"11001100",	-- ##..##..
		1189 =>	"11001100",	-- ##..##..
		1190 =>	"01111000",	-- .####...
		1191 =>	"00000000",	-- ........

		-- char 0x95='\x95
		1192 =>	"01100000",	-- .##.....
		1193 =>	"00110000",	-- ..##....
		1194 =>	"00000000",	-- ........
		1195 =>	"01111000",	-- .####...
		1196 =>	"11001100",	-- ##..##..
		1197 =>	"11001100",	-- ##..##..
		1198 =>	"01111000",	-- .####...
		1199 =>	"00000000",	-- ........

		-- char 0x96='\x96
		1200 =>	"01111000",	-- .####...
		1201 =>	"11001100",	-- ##..##..
		1202 =>	"00000000",	-- ........
		1203 =>	"11001100",	-- ##..##..
		1204 =>	"11001100",	-- ##..##..
		1205 =>	"11001100",	-- ##..##..
		1206 =>	"01111110",	-- .######.
		1207 =>	"00000000",	-- ........

		-- char 0x97='\x97
		1208 =>	"01100000",	-- .##.....
		1209 =>	"00110000",	-- ..##....
		1210 =>	"00000000",	-- ........
		1211 =>	"11001100",	-- ##..##..
		1212 =>	"11001100",	-- ##..##..
		1213 =>	"11001100",	-- ##..##..
		1214 =>	"01111110",	-- .######.
		1215 =>	"00000000",	-- ........

		-- char 0x98='\x98
		1216 =>	"00000000",	-- ........
		1217 =>	"11001100",	-- ##..##..
		1218 =>	"00000000",	-- ........
		1219 =>	"11001100",	-- ##..##..
		1220 =>	"11001100",	-- ##..##..
		1221 =>	"11111100",	-- ######..
		1222 =>	"00001100",	-- ....##..
		1223 =>	"11111000",	-- #####...

		-- char 0x99='\x99
		1224 =>	"11000110",	-- ##...##.
		1225 =>	"00000000",	-- ........
		1226 =>	"01111100",	-- .#####..
		1227 =>	"11000110",	-- ##...##.
		1228 =>	"11000110",	-- ##...##.
		1229 =>	"11000110",	-- ##...##.
		1230 =>	"01111100",	-- .#####..
		1231 =>	"00000000",	-- ........

		-- char 0x9a='\x9a
		1232 =>	"11001100",	-- ##..##..
		1233 =>	"00000000",	-- ........
		1234 =>	"11001100",	-- ##..##..
		1235 =>	"11001100",	-- ##..##..
		1236 =>	"11001100",	-- ##..##..
		1237 =>	"11001100",	-- ##..##..
		1238 =>	"01111000",	-- .####...
		1239 =>	"00000000",	-- ........

		-- char 0x9b='\x9b
		1240 =>	"00011000",	-- ...##...
		1241 =>	"00011000",	-- ...##...
		1242 =>	"01111110",	-- .######.
		1243 =>	"11000000",	-- ##......
		1244 =>	"11000000",	-- ##......
		1245 =>	"01111110",	-- .######.
		1246 =>	"00011000",	-- ...##...
		1247 =>	"00011000",	-- ...##...

		-- char 0x9c='\x9c
		1248 =>	"00111000",	-- ..###...
		1249 =>	"01101100",	-- .##.##..
		1250 =>	"01100100",	-- .##..#..
		1251 =>	"11110000",	-- ####....
		1252 =>	"01100000",	-- .##.....
		1253 =>	"11100110",	-- ###..##.
		1254 =>	"11111100",	-- ######..
		1255 =>	"00000000",	-- ........

		-- char 0x9d='\x9d
		1256 =>	"11001100",	-- ##..##..
		1257 =>	"11001100",	-- ##..##..
		1258 =>	"01111000",	-- .####...
		1259 =>	"11111100",	-- ######..
		1260 =>	"00110000",	-- ..##....
		1261 =>	"11111100",	-- ######..
		1262 =>	"00110000",	-- ..##....
		1263 =>	"00110000",	-- ..##....

		-- char 0x9e='\x9e
		1264 =>	"00000000",	-- ........
		1265 =>	"00000000",	-- ........
		1266 =>	"11001100",	-- ##..##..
		1267 =>	"01111000",	-- .####...
		1268 =>	"00110000",	-- ..##....
		1269 =>	"01111000",	-- .####...
		1270 =>	"11001100",	-- ##..##..
		1271 =>	"00000000",	-- ........

		-- char 0x9f='\x9f
		1272 =>	"00001110",	-- ....###.
		1273 =>	"00011011",	-- ...##.##
		1274 =>	"00011000",	-- ...##...
		1275 =>	"01111110",	-- .######.
		1276 =>	"00011000",	-- ...##...
		1277 =>	"00011000",	-- ...##...
		1278 =>	"11011000",	-- ##.##...
		1279 =>	"01110000",	-- .###....

		-- char 0xa0='\xa0
		1280 =>	"00011000",	-- ...##...
		1281 =>	"00110000",	-- ..##....
		1282 =>	"01111000",	-- .####...
		1283 =>	"00001100",	-- ....##..
		1284 =>	"01111100",	-- .#####..
		1285 =>	"11001100",	-- ##..##..
		1286 =>	"01111110",	-- .######.
		1287 =>	"00000000",	-- ........

		-- char 0xa1='\xa1
		1288 =>	"00011000",	-- ...##...
		1289 =>	"00110000",	-- ..##....
		1290 =>	"01110000",	-- .###....
		1291 =>	"00110000",	-- ..##....
		1292 =>	"00110000",	-- ..##....
		1293 =>	"00110000",	-- ..##....
		1294 =>	"01111000",	-- .####...
		1295 =>	"00000000",	-- ........

		-- char 0xa2='\xa2
		1296 =>	"00001100",	-- ....##..
		1297 =>	"00011000",	-- ...##...
		1298 =>	"00000000",	-- ........
		1299 =>	"01111000",	-- .####...
		1300 =>	"11001100",	-- ##..##..
		1301 =>	"11001100",	-- ##..##..
		1302 =>	"01111000",	-- .####...
		1303 =>	"00000000",	-- ........

		-- char 0xa3='\xa3
		1304 =>	"00001100",	-- ....##..
		1305 =>	"00011000",	-- ...##...
		1306 =>	"00000000",	-- ........
		1307 =>	"11001100",	-- ##..##..
		1308 =>	"11001100",	-- ##..##..
		1309 =>	"11001100",	-- ##..##..
		1310 =>	"01111110",	-- .######.
		1311 =>	"00000000",	-- ........

		-- char 0xa4='\xa4
		1312 =>	"01110110",	-- .###.##.
		1313 =>	"11011100",	-- ##.###..
		1314 =>	"00000000",	-- ........
		1315 =>	"11111000",	-- #####...
		1316 =>	"11001100",	-- ##..##..
		1317 =>	"11001100",	-- ##..##..
		1318 =>	"11001100",	-- ##..##..
		1319 =>	"00000000",	-- ........

		-- char 0xa5='\xa5
		1320 =>	"01110110",	-- .###.##.
		1321 =>	"11011100",	-- ##.###..
		1322 =>	"00000000",	-- ........
		1323 =>	"11101100",	-- ###.##..
		1324 =>	"11111100",	-- ######..
		1325 =>	"11011100",	-- ##.###..
		1326 =>	"11001100",	-- ##..##..
		1327 =>	"00000000",	-- ........

		-- char 0xa6='\xa6
		1328 =>	"00111100",	-- ..####..
		1329 =>	"01101100",	-- .##.##..
		1330 =>	"01101100",	-- .##.##..
		1331 =>	"00111110",	-- ..#####.
		1332 =>	"00000000",	-- ........
		1333 =>	"01111110",	-- .######.
		1334 =>	"00000000",	-- ........
		1335 =>	"00000000",	-- ........

		-- char 0xa7='\xa7
		1336 =>	"00111100",	-- ..####..
		1337 =>	"01100110",	-- .##..##.
		1338 =>	"01100110",	-- .##..##.
		1339 =>	"00111100",	-- ..####..
		1340 =>	"00000000",	-- ........
		1341 =>	"01111110",	-- .######.
		1342 =>	"00000000",	-- ........
		1343 =>	"00000000",	-- ........

		-- char 0xa8='\xa8
		1344 =>	"00110000",	-- ..##....
		1345 =>	"00000000",	-- ........
		1346 =>	"00110000",	-- ..##....
		1347 =>	"01100000",	-- .##.....
		1348 =>	"11000000",	-- ##......
		1349 =>	"11001100",	-- ##..##..
		1350 =>	"01111000",	-- .####...
		1351 =>	"00000000",	-- ........

		-- char 0xa9='\xa9
		1352 =>	"00000000",	-- ........
		1353 =>	"00000000",	-- ........
		1354 =>	"00000000",	-- ........
		1355 =>	"11111100",	-- ######..
		1356 =>	"11000000",	-- ##......
		1357 =>	"11000000",	-- ##......
		1358 =>	"00000000",	-- ........
		1359 =>	"00000000",	-- ........

		-- char 0xaa='\xaa
		1360 =>	"00000000",	-- ........
		1361 =>	"00000000",	-- ........
		1362 =>	"00000000",	-- ........
		1363 =>	"11111100",	-- ######..
		1364 =>	"00001100",	-- ....##..
		1365 =>	"00001100",	-- ....##..
		1366 =>	"00000000",	-- ........
		1367 =>	"00000000",	-- ........

		-- char 0xab='\xab
		1368 =>	"11000011",	-- ##....##
		1369 =>	"11000110",	-- ##...##.
		1370 =>	"11001100",	-- ##..##..
		1371 =>	"11011110",	-- ##.####.
		1372 =>	"00110011",	-- ..##..##
		1373 =>	"01100110",	-- .##..##.
		1374 =>	"11001100",	-- ##..##..
		1375 =>	"00001111",	-- ....####

		-- char 0xac='\xac
		1376 =>	"11000011",	-- ##....##
		1377 =>	"11000110",	-- ##...##.
		1378 =>	"11001100",	-- ##..##..
		1379 =>	"11011011",	-- ##.##.##
		1380 =>	"00110111",	-- ..##.###
		1381 =>	"01101111",	-- .##.####
		1382 =>	"11001111",	-- ##..####
		1383 =>	"00000011",	-- ......##

		-- char 0xad='\xad
		1384 =>	"00000000",	-- ........
		1385 =>	"00011000",	-- ...##...
		1386 =>	"00000000",	-- ........
		1387 =>	"00011000",	-- ...##...
		1388 =>	"00011000",	-- ...##...
		1389 =>	"00111100",	-- ..####..
		1390 =>	"00111100",	-- ..####..
		1391 =>	"00011000",	-- ...##...

		-- char 0xae='\xae
		1392 =>	"00000000",	-- ........
		1393 =>	"00110011",	-- ..##..##
		1394 =>	"01100110",	-- .##..##.
		1395 =>	"11001100",	-- ##..##..
		1396 =>	"01100110",	-- .##..##.
		1397 =>	"00110011",	-- ..##..##
		1398 =>	"00000000",	-- ........
		1399 =>	"00000000",	-- ........

		-- char 0xaf='\xaf
		1400 =>	"00000000",	-- ........
		1401 =>	"11001100",	-- ##..##..
		1402 =>	"01100110",	-- .##..##.
		1403 =>	"00110011",	-- ..##..##
		1404 =>	"01100110",	-- .##..##.
		1405 =>	"11001100",	-- ##..##..
		1406 =>	"00000000",	-- ........
		1407 =>	"00000000",	-- ........

		-- char 0xb0='\xb0
		1408 =>	"00100010",	-- ..#...#.
		1409 =>	"10001000",	-- #...#...
		1410 =>	"00100010",	-- ..#...#.
		1411 =>	"10001000",	-- #...#...
		1412 =>	"00100010",	-- ..#...#.
		1413 =>	"10001000",	-- #...#...
		1414 =>	"00100010",	-- ..#...#.
		1415 =>	"10001000",	-- #...#...

		-- char 0xb1='\xb1
		1416 =>	"01010101",	-- .#.#.#.#
		1417 =>	"10101010",	-- #.#.#.#.
		1418 =>	"01010101",	-- .#.#.#.#
		1419 =>	"10101010",	-- #.#.#.#.
		1420 =>	"01010101",	-- .#.#.#.#
		1421 =>	"10101010",	-- #.#.#.#.
		1422 =>	"01010101",	-- .#.#.#.#
		1423 =>	"10101010",	-- #.#.#.#.

		-- char 0xb2='\xb2
		1424 =>	"11011101",	-- ##.###.#
		1425 =>	"01110111",	-- .###.###
		1426 =>	"11011101",	-- ##.###.#
		1427 =>	"01110111",	-- .###.###
		1428 =>	"11011101",	-- ##.###.#
		1429 =>	"01110111",	-- .###.###
		1430 =>	"11011101",	-- ##.###.#
		1431 =>	"01110111",	-- .###.###

		-- char 0xb3='\xb3
		1432 =>	"00011000",	-- ...##...
		1433 =>	"00011000",	-- ...##...
		1434 =>	"00011000",	-- ...##...
		1435 =>	"00011000",	-- ...##...
		1436 =>	"00011000",	-- ...##...
		1437 =>	"00011000",	-- ...##...
		1438 =>	"00011000",	-- ...##...
		1439 =>	"00011000",	-- ...##...

		-- char 0xb4='\xb4
		1440 =>	"00011000",	-- ...##...
		1441 =>	"00011000",	-- ...##...
		1442 =>	"00011000",	-- ...##...
		1443 =>	"11111000",	-- #####...
		1444 =>	"11111000",	-- #####...
		1445 =>	"00011000",	-- ...##...
		1446 =>	"00011000",	-- ...##...
		1447 =>	"00011000",	-- ...##...

		-- char 0xb5='\xb5
		1448 =>	"00011000",	-- ...##...
		1449 =>	"11111000",	-- #####...
		1450 =>	"11111000",	-- #####...
		1451 =>	"00011000",	-- ...##...
		1452 =>	"00011000",	-- ...##...
		1453 =>	"11111000",	-- #####...
		1454 =>	"11111000",	-- #####...
		1455 =>	"00011000",	-- ...##...

		-- char 0xb6='\xb6
		1456 =>	"01100110",	-- .##..##.
		1457 =>	"01100110",	-- .##..##.
		1458 =>	"01100110",	-- .##..##.
		1459 =>	"11100110",	-- ###..##.
		1460 =>	"11100110",	-- ###..##.
		1461 =>	"01100110",	-- .##..##.
		1462 =>	"01100110",	-- .##..##.
		1463 =>	"01100110",	-- .##..##.

		-- char 0xb7='\xb7
		1464 =>	"00000000",	-- ........
		1465 =>	"00000000",	-- ........
		1466 =>	"00000000",	-- ........
		1467 =>	"11111110",	-- #######.
		1468 =>	"11111110",	-- #######.
		1469 =>	"01100110",	-- .##..##.
		1470 =>	"01100110",	-- .##..##.
		1471 =>	"01100110",	-- .##..##.

		-- char 0xb8='\xb8
		1472 =>	"00000000",	-- ........
		1473 =>	"11111000",	-- #####...
		1474 =>	"11111000",	-- #####...
		1475 =>	"00011000",	-- ...##...
		1476 =>	"00011000",	-- ...##...
		1477 =>	"11111000",	-- #####...
		1478 =>	"11111000",	-- #####...
		1479 =>	"00011000",	-- ...##...

		-- char 0xb9='\xb9
		1480 =>	"01100110",	-- .##..##.
		1481 =>	"11100110",	-- ###..##.
		1482 =>	"11100110",	-- ###..##.
		1483 =>	"00000110",	-- .....##.
		1484 =>	"00000110",	-- .....##.
		1485 =>	"11100110",	-- ###..##.
		1486 =>	"11100110",	-- ###..##.
		1487 =>	"01100110",	-- .##..##.

		-- char 0xba='\xba
		1488 =>	"01100110",	-- .##..##.
		1489 =>	"01100110",	-- .##..##.
		1490 =>	"01100110",	-- .##..##.
		1491 =>	"01100110",	-- .##..##.
		1492 =>	"01100110",	-- .##..##.
		1493 =>	"01100110",	-- .##..##.
		1494 =>	"01100110",	-- .##..##.
		1495 =>	"01100110",	-- .##..##.

		-- char 0xbb='\xbb
		1496 =>	"00000000",	-- ........
		1497 =>	"11111110",	-- #######.
		1498 =>	"11111110",	-- #######.
		1499 =>	"00000110",	-- .....##.
		1500 =>	"00000110",	-- .....##.
		1501 =>	"11100110",	-- ###..##.
		1502 =>	"11100110",	-- ###..##.
		1503 =>	"01100110",	-- .##..##.

		-- char 0xbc='\xbc
		1504 =>	"01100110",	-- .##..##.
		1505 =>	"11100110",	-- ###..##.
		1506 =>	"11100110",	-- ###..##.
		1507 =>	"00000110",	-- .....##.
		1508 =>	"00000110",	-- .....##.
		1509 =>	"11111110",	-- #######.
		1510 =>	"11111110",	-- #######.
		1511 =>	"00000000",	-- ........

		-- char 0xbd='\xbd
		1512 =>	"01100110",	-- .##..##.
		1513 =>	"01100110",	-- .##..##.
		1514 =>	"01100110",	-- .##..##.
		1515 =>	"01100110",	-- .##..##.
		1516 =>	"11111110",	-- #######.
		1517 =>	"11111110",	-- #######.
		1518 =>	"00000000",	-- ........
		1519 =>	"00000000",	-- ........

		-- char 0xbe='\xbe
		1520 =>	"00011000",	-- ...##...
		1521 =>	"11111000",	-- #####...
		1522 =>	"11111000",	-- #####...
		1523 =>	"00011000",	-- ...##...
		1524 =>	"00011000",	-- ...##...
		1525 =>	"11111000",	-- #####...
		1526 =>	"11111000",	-- #####...
		1527 =>	"00000000",	-- ........

		-- char 0xbf='\xbf
		1528 =>	"00000000",	-- ........
		1529 =>	"00000000",	-- ........
		1530 =>	"00000000",	-- ........
		1531 =>	"11111000",	-- #####...
		1532 =>	"11111000",	-- #####...
		1533 =>	"00011000",	-- ...##...
		1534 =>	"00011000",	-- ...##...
		1535 =>	"00011000",	-- ...##...

		-- char 0xc0='\xc0
		1536 =>	"00011000",	-- ...##...
		1537 =>	"00011000",	-- ...##...
		1538 =>	"00011000",	-- ...##...
		1539 =>	"00011111",	-- ...#####
		1540 =>	"00011111",	-- ...#####
		1541 =>	"00000000",	-- ........
		1542 =>	"00000000",	-- ........
		1543 =>	"00000000",	-- ........

		-- char 0xc1='\xc1
		1544 =>	"00011000",	-- ...##...
		1545 =>	"00011000",	-- ...##...
		1546 =>	"00011000",	-- ...##...
		1547 =>	"11111111",	-- ########
		1548 =>	"11111111",	-- ########
		1549 =>	"00000000",	-- ........
		1550 =>	"00000000",	-- ........
		1551 =>	"00000000",	-- ........

		-- char 0xc2='\xc2
		1552 =>	"00000000",	-- ........
		1553 =>	"00000000",	-- ........
		1554 =>	"00000000",	-- ........
		1555 =>	"11111111",	-- ########
		1556 =>	"11111111",	-- ########
		1557 =>	"00011000",	-- ...##...
		1558 =>	"00011000",	-- ...##...
		1559 =>	"00011000",	-- ...##...

		-- char 0xc3='\xc3
		1560 =>	"00011000",	-- ...##...
		1561 =>	"00011000",	-- ...##...
		1562 =>	"00011000",	-- ...##...
		1563 =>	"00011111",	-- ...#####
		1564 =>	"00011111",	-- ...#####
		1565 =>	"00011000",	-- ...##...
		1566 =>	"00011000",	-- ...##...
		1567 =>	"00011000",	-- ...##...

		-- char 0xc4='\xc4
		1568 =>	"00000000",	-- ........
		1569 =>	"00000000",	-- ........
		1570 =>	"00000000",	-- ........
		1571 =>	"11111111",	-- ########
		1572 =>	"11111111",	-- ########
		1573 =>	"00000000",	-- ........
		1574 =>	"00000000",	-- ........
		1575 =>	"00000000",	-- ........

		-- char 0xc5='\xc5
		1576 =>	"00011000",	-- ...##...
		1577 =>	"00011000",	-- ...##...
		1578 =>	"00011000",	-- ...##...
		1579 =>	"11111111",	-- ########
		1580 =>	"11111111",	-- ########
		1581 =>	"00011000",	-- ...##...
		1582 =>	"00011000",	-- ...##...
		1583 =>	"00011000",	-- ...##...

		-- char 0xc6='\xc6
		1584 =>	"00011000",	-- ...##...
		1585 =>	"00011111",	-- ...#####
		1586 =>	"00011111",	-- ...#####
		1587 =>	"00011000",	-- ...##...
		1588 =>	"00011000",	-- ...##...
		1589 =>	"00011111",	-- ...#####
		1590 =>	"00011111",	-- ...#####
		1591 =>	"00011000",	-- ...##...

		-- char 0xc7='\xc7
		1592 =>	"01100110",	-- .##..##.
		1593 =>	"01100110",	-- .##..##.
		1594 =>	"01100110",	-- .##..##.
		1595 =>	"01100111",	-- .##..###
		1596 =>	"01100111",	-- .##..###
		1597 =>	"01100110",	-- .##..##.
		1598 =>	"01100110",	-- .##..##.
		1599 =>	"01100110",	-- .##..##.

		-- char 0xc8='\xc8
		1600 =>	"01100110",	-- .##..##.
		1601 =>	"01100111",	-- .##..###
		1602 =>	"01100111",	-- .##..###
		1603 =>	"01100000",	-- .##.....
		1604 =>	"01100000",	-- .##.....
		1605 =>	"01111111",	-- .#######
		1606 =>	"01111111",	-- .#######
		1607 =>	"00000000",	-- ........

		-- char 0xc9='\xc9
		1608 =>	"00000000",	-- ........
		1609 =>	"01111111",	-- .#######
		1610 =>	"01111111",	-- .#######
		1611 =>	"01100000",	-- .##.....
		1612 =>	"01100000",	-- .##.....
		1613 =>	"01100111",	-- .##..###
		1614 =>	"01100111",	-- .##..###
		1615 =>	"01100110",	-- .##..##.

		-- char 0xca='\xca
		1616 =>	"01100110",	-- .##..##.
		1617 =>	"11100111",	-- ###..###
		1618 =>	"11100111",	-- ###..###
		1619 =>	"00000000",	-- ........
		1620 =>	"00000000",	-- ........
		1621 =>	"11111111",	-- ########
		1622 =>	"11111111",	-- ########
		1623 =>	"00000000",	-- ........

		-- char 0xcb='\xcb
		1624 =>	"00000000",	-- ........
		1625 =>	"11111111",	-- ########
		1626 =>	"11111111",	-- ########
		1627 =>	"00000000",	-- ........
		1628 =>	"00000000",	-- ........
		1629 =>	"11100111",	-- ###..###
		1630 =>	"11100111",	-- ###..###
		1631 =>	"01100110",	-- .##..##.

		-- char 0xcc='\xcc
		1632 =>	"01100110",	-- .##..##.
		1633 =>	"01100111",	-- .##..###
		1634 =>	"01100111",	-- .##..###
		1635 =>	"01100000",	-- .##.....
		1636 =>	"01100000",	-- .##.....
		1637 =>	"01100111",	-- .##..###
		1638 =>	"01100111",	-- .##..###
		1639 =>	"01100110",	-- .##..##.

		-- char 0xcd='\xcd
		1640 =>	"00000000",	-- ........
		1641 =>	"11111111",	-- ########
		1642 =>	"11111111",	-- ########
		1643 =>	"00000000",	-- ........
		1644 =>	"00000000",	-- ........
		1645 =>	"11111111",	-- ########
		1646 =>	"11111111",	-- ########
		1647 =>	"00000000",	-- ........

		-- char 0xce='\xce
		1648 =>	"01100110",	-- .##..##.
		1649 =>	"11100111",	-- ###..###
		1650 =>	"11100111",	-- ###..###
		1651 =>	"00000000",	-- ........
		1652 =>	"00000000",	-- ........
		1653 =>	"11100111",	-- ###..###
		1654 =>	"11100111",	-- ###..###
		1655 =>	"01100110",	-- .##..##.

		-- char 0xcf='\xcf
		1656 =>	"00011000",	-- ...##...
		1657 =>	"11111111",	-- ########
		1658 =>	"11111111",	-- ########
		1659 =>	"00000000",	-- ........
		1660 =>	"00000000",	-- ........
		1661 =>	"11111111",	-- ########
		1662 =>	"11111111",	-- ########
		1663 =>	"00000000",	-- ........

		-- char 0xd0='\xd0
		1664 =>	"01100110",	-- .##..##.
		1665 =>	"01100110",	-- .##..##.
		1666 =>	"01100110",	-- .##..##.
		1667 =>	"11111111",	-- ########
		1668 =>	"11111111",	-- ########
		1669 =>	"00000000",	-- ........
		1670 =>	"00000000",	-- ........
		1671 =>	"00000000",	-- ........

		-- char 0xd1='\xd1
		1672 =>	"00000000",	-- ........
		1673 =>	"11111111",	-- ########
		1674 =>	"11111111",	-- ########
		1675 =>	"00000000",	-- ........
		1676 =>	"00000000",	-- ........
		1677 =>	"11111111",	-- ########
		1678 =>	"11111111",	-- ########
		1679 =>	"00011000",	-- ...##...

		-- char 0xd2='\xd2
		1680 =>	"00000000",	-- ........
		1681 =>	"00000000",	-- ........
		1682 =>	"00000000",	-- ........
		1683 =>	"00000000",	-- ........
		1684 =>	"00000000",	-- ........
		1685 =>	"11111111",	-- ########
		1686 =>	"11111111",	-- ########
		1687 =>	"01100110",	-- .##..##.

		-- char 0xd3='\xd3
		1688 =>	"01100110",	-- .##..##.
		1689 =>	"01100110",	-- .##..##.
		1690 =>	"01100110",	-- .##..##.
		1691 =>	"01111111",	-- .#######
		1692 =>	"01111111",	-- .#######
		1693 =>	"00000000",	-- ........
		1694 =>	"00000000",	-- ........
		1695 =>	"00000000",	-- ........

		-- char 0xd4='\xd4
		1696 =>	"00011000",	-- ...##...
		1697 =>	"00011111",	-- ...#####
		1698 =>	"00011111",	-- ...#####
		1699 =>	"00011000",	-- ...##...
		1700 =>	"00011000",	-- ...##...
		1701 =>	"00011111",	-- ...#####
		1702 =>	"00011111",	-- ...#####
		1703 =>	"00000000",	-- ........

		-- char 0xd5='\xd5
		1704 =>	"00000000",	-- ........
		1705 =>	"00011111",	-- ...#####
		1706 =>	"00011111",	-- ...#####
		1707 =>	"00011000",	-- ...##...
		1708 =>	"00011000",	-- ...##...
		1709 =>	"00011111",	-- ...#####
		1710 =>	"00011111",	-- ...#####
		1711 =>	"00011000",	-- ...##...

		-- char 0xd6='\xd6
		1712 =>	"00000000",	-- ........
		1713 =>	"00000000",	-- ........
		1714 =>	"00000000",	-- ........
		1715 =>	"01111111",	-- .#######
		1716 =>	"01111111",	-- .#######
		1717 =>	"01100110",	-- .##..##.
		1718 =>	"01100110",	-- .##..##.
		1719 =>	"01100110",	-- .##..##.

		-- char 0xd7='\xd7
		1720 =>	"01100110",	-- .##..##.
		1721 =>	"01100110",	-- .##..##.
		1722 =>	"01100110",	-- .##..##.
		1723 =>	"11111111",	-- ########
		1724 =>	"11111111",	-- ########
		1725 =>	"01100110",	-- .##..##.
		1726 =>	"01100110",	-- .##..##.
		1727 =>	"01100110",	-- .##..##.

		-- char 0xd8='\xd8
		1728 =>	"00011000",	-- ...##...
		1729 =>	"11111111",	-- ########
		1730 =>	"11111111",	-- ########
		1731 =>	"00011000",	-- ...##...
		1732 =>	"00011000",	-- ...##...
		1733 =>	"11111111",	-- ########
		1734 =>	"11111111",	-- ########
		1735 =>	"00011000",	-- ...##...

		-- char 0xd9='\xd9
		1736 =>	"00011000",	-- ...##...
		1737 =>	"00011000",	-- ...##...
		1738 =>	"00011000",	-- ...##...
		1739 =>	"11111000",	-- #####...
		1740 =>	"11111000",	-- #####...
		1741 =>	"00000000",	-- ........
		1742 =>	"00000000",	-- ........
		1743 =>	"00000000",	-- ........

		-- char 0xda='\xda
		1744 =>	"00000000",	-- ........
		1745 =>	"00000000",	-- ........
		1746 =>	"00000000",	-- ........
		1747 =>	"00011111",	-- ...#####
		1748 =>	"00011111",	-- ...#####
		1749 =>	"00011000",	-- ...##...
		1750 =>	"00011000",	-- ...##...
		1751 =>	"00011000",	-- ...##...

		-- char 0xdb='\xdb
		1752 =>	"11111111",	-- ########
		1753 =>	"11111111",	-- ########
		1754 =>	"11111111",	-- ########
		1755 =>	"11111111",	-- ########
		1756 =>	"11111111",	-- ########
		1757 =>	"11111111",	-- ########
		1758 =>	"11111111",	-- ########
		1759 =>	"11111111",	-- ########

		-- char 0xdc='\xdc
		1760 =>	"00000000",	-- ........
		1761 =>	"00000000",	-- ........
		1762 =>	"00000000",	-- ........
		1763 =>	"00000000",	-- ........
		1764 =>	"11111111",	-- ########
		1765 =>	"11111111",	-- ########
		1766 =>	"11111111",	-- ########
		1767 =>	"11111111",	-- ########

		-- char 0xdd='\xdd
		1768 =>	"11110000",	-- ####....
		1769 =>	"11110000",	-- ####....
		1770 =>	"11110000",	-- ####....
		1771 =>	"11110000",	-- ####....
		1772 =>	"11110000",	-- ####....
		1773 =>	"11110000",	-- ####....
		1774 =>	"11110000",	-- ####....
		1775 =>	"11110000",	-- ####....

		-- char 0xde='\xde
		1776 =>	"00001111",	-- ....####
		1777 =>	"00001111",	-- ....####
		1778 =>	"00001111",	-- ....####
		1779 =>	"00001111",	-- ....####
		1780 =>	"00001111",	-- ....####
		1781 =>	"00001111",	-- ....####
		1782 =>	"00001111",	-- ....####
		1783 =>	"00001111",	-- ....####

		-- char 0xdf='\xdf
		1784 =>	"11111111",	-- ########
		1785 =>	"11111111",	-- ########
		1786 =>	"11111111",	-- ########
		1787 =>	"11111111",	-- ########
		1788 =>	"00000000",	-- ........
		1789 =>	"00000000",	-- ........
		1790 =>	"00000000",	-- ........
		1791 =>	"00000000",	-- ........

		-- char 0xe0='\xe0
		1792 =>	"00000000",	-- ........
		1793 =>	"00000000",	-- ........
		1794 =>	"01110110",	-- .###.##.
		1795 =>	"11011100",	-- ##.###..
		1796 =>	"11001000",	-- ##..#...
		1797 =>	"11011100",	-- ##.###..
		1798 =>	"01110110",	-- .###.##.
		1799 =>	"00000000",	-- ........

		-- char 0xe1='\xe1
		1800 =>	"00000000",	-- ........
		1801 =>	"01111000",	-- .####...
		1802 =>	"11001100",	-- ##..##..
		1803 =>	"11111000",	-- #####...
		1804 =>	"11001100",	-- ##..##..
		1805 =>	"11111000",	-- #####...
		1806 =>	"11000000",	-- ##......
		1807 =>	"11000000",	-- ##......

		-- char 0xe2='\xe2
		1808 =>	"00000000",	-- ........
		1809 =>	"11111100",	-- ######..
		1810 =>	"11001100",	-- ##..##..
		1811 =>	"11000000",	-- ##......
		1812 =>	"11000000",	-- ##......
		1813 =>	"11000000",	-- ##......
		1814 =>	"11000000",	-- ##......
		1815 =>	"00000000",	-- ........

		-- char 0xe3='\xe3
		1816 =>	"00000000",	-- ........
		1817 =>	"11111110",	-- #######.
		1818 =>	"01101100",	-- .##.##..
		1819 =>	"01101100",	-- .##.##..
		1820 =>	"01101100",	-- .##.##..
		1821 =>	"01101100",	-- .##.##..
		1822 =>	"01101100",	-- .##.##..
		1823 =>	"00000000",	-- ........

		-- char 0xe4='\xe4
		1824 =>	"11111100",	-- ######..
		1825 =>	"11001100",	-- ##..##..
		1826 =>	"01100000",	-- .##.....
		1827 =>	"00110000",	-- ..##....
		1828 =>	"01100000",	-- .##.....
		1829 =>	"11001100",	-- ##..##..
		1830 =>	"11111100",	-- ######..
		1831 =>	"00000000",	-- ........

		-- char 0xe5='\xe5
		1832 =>	"00000000",	-- ........
		1833 =>	"00000000",	-- ........
		1834 =>	"01111110",	-- .######.
		1835 =>	"11011000",	-- ##.##...
		1836 =>	"11011000",	-- ##.##...
		1837 =>	"11011000",	-- ##.##...
		1838 =>	"01110000",	-- .###....
		1839 =>	"00000000",	-- ........

		-- char 0xe6='\xe6
		1840 =>	"00000000",	-- ........
		1841 =>	"01100110",	-- .##..##.
		1842 =>	"01100110",	-- .##..##.
		1843 =>	"01100110",	-- .##..##.
		1844 =>	"01100110",	-- .##..##.
		1845 =>	"01111100",	-- .#####..
		1846 =>	"01100000",	-- .##.....
		1847 =>	"11000000",	-- ##......

		-- char 0xe7='\xe7
		1848 =>	"00000000",	-- ........
		1849 =>	"01110110",	-- .###.##.
		1850 =>	"11011100",	-- ##.###..
		1851 =>	"00011000",	-- ...##...
		1852 =>	"00011000",	-- ...##...
		1853 =>	"00011000",	-- ...##...
		1854 =>	"00011000",	-- ...##...
		1855 =>	"00000000",	-- ........

		-- char 0xe8='\xe8
		1856 =>	"11111100",	-- ######..
		1857 =>	"00110000",	-- ..##....
		1858 =>	"01111000",	-- .####...
		1859 =>	"11001100",	-- ##..##..
		1860 =>	"11001100",	-- ##..##..
		1861 =>	"01111000",	-- .####...
		1862 =>	"00110000",	-- ..##....
		1863 =>	"11111100",	-- ######..

		-- char 0xe9='\xe9
		1864 =>	"00111000",	-- ..###...
		1865 =>	"01101100",	-- .##.##..
		1866 =>	"11000110",	-- ##...##.
		1867 =>	"11111110",	-- #######.
		1868 =>	"11000110",	-- ##...##.
		1869 =>	"01101100",	-- .##.##..
		1870 =>	"00111000",	-- ..###...
		1871 =>	"00000000",	-- ........

		-- char 0xea='\xea
		1872 =>	"00111000",	-- ..###...
		1873 =>	"01101100",	-- .##.##..
		1874 =>	"11000110",	-- ##...##.
		1875 =>	"11000110",	-- ##...##.
		1876 =>	"01101100",	-- .##.##..
		1877 =>	"01101100",	-- .##.##..
		1878 =>	"11101110",	-- ###.###.
		1879 =>	"00000000",	-- ........

		-- char 0xeb='\xeb
		1880 =>	"00011100",	-- ...###..
		1881 =>	"00110000",	-- ..##....
		1882 =>	"00011000",	-- ...##...
		1883 =>	"01111100",	-- .#####..
		1884 =>	"11001100",	-- ##..##..
		1885 =>	"11001100",	-- ##..##..
		1886 =>	"01111000",	-- .####...
		1887 =>	"00000000",	-- ........

		-- char 0xec='\xec
		1888 =>	"00000000",	-- ........
		1889 =>	"00000000",	-- ........
		1890 =>	"01111110",	-- .######.
		1891 =>	"11011011",	-- ##.##.##
		1892 =>	"11011011",	-- ##.##.##
		1893 =>	"01111110",	-- .######.
		1894 =>	"00000000",	-- ........
		1895 =>	"00000000",	-- ........

		-- char 0xed='\xed
		1896 =>	"00000110",	-- .....##.
		1897 =>	"00001100",	-- ....##..
		1898 =>	"01111110",	-- .######.
		1899 =>	"11011011",	-- ##.##.##
		1900 =>	"11011011",	-- ##.##.##
		1901 =>	"01111110",	-- .######.
		1902 =>	"01100000",	-- .##.....
		1903 =>	"11000000",	-- ##......

		-- char 0xee='\xee
		1904 =>	"00111000",	-- ..###...
		1905 =>	"01100000",	-- .##.....
		1906 =>	"11000000",	-- ##......
		1907 =>	"11111000",	-- #####...
		1908 =>	"11000000",	-- ##......
		1909 =>	"01100000",	-- .##.....
		1910 =>	"00111000",	-- ..###...
		1911 =>	"00000000",	-- ........

		-- char 0xef='\xef
		1912 =>	"01111000",	-- .####...
		1913 =>	"11001100",	-- ##..##..
		1914 =>	"11001100",	-- ##..##..
		1915 =>	"11001100",	-- ##..##..
		1916 =>	"11001100",	-- ##..##..
		1917 =>	"11001100",	-- ##..##..
		1918 =>	"11001100",	-- ##..##..
		1919 =>	"00000000",	-- ........

		-- char 0xf0='\xf0
		1920 =>	"00000000",	-- ........
		1921 =>	"11111100",	-- ######..
		1922 =>	"00000000",	-- ........
		1923 =>	"11111100",	-- ######..
		1924 =>	"00000000",	-- ........
		1925 =>	"11111100",	-- ######..
		1926 =>	"00000000",	-- ........
		1927 =>	"00000000",	-- ........

		-- char 0xf1='\xf1
		1928 =>	"00110000",	-- ..##....
		1929 =>	"00110000",	-- ..##....
		1930 =>	"11111100",	-- ######..
		1931 =>	"00110000",	-- ..##....
		1932 =>	"00110000",	-- ..##....
		1933 =>	"00000000",	-- ........
		1934 =>	"11111100",	-- ######..
		1935 =>	"00000000",	-- ........

		-- char 0xf2='\xf2
		1936 =>	"01100000",	-- .##.....
		1937 =>	"00110000",	-- ..##....
		1938 =>	"00011000",	-- ...##...
		1939 =>	"00110000",	-- ..##....
		1940 =>	"01100000",	-- .##.....
		1941 =>	"00000000",	-- ........
		1942 =>	"11111100",	-- ######..
		1943 =>	"00000000",	-- ........

		-- char 0xf3='\xf3
		1944 =>	"00011000",	-- ...##...
		1945 =>	"00110000",	-- ..##....
		1946 =>	"01100000",	-- .##.....
		1947 =>	"00110000",	-- ..##....
		1948 =>	"00011000",	-- ...##...
		1949 =>	"00000000",	-- ........
		1950 =>	"11111100",	-- ######..
		1951 =>	"00000000",	-- ........

		-- char 0xf4='\xf4
		1952 =>	"00001110",	-- ....###.
		1953 =>	"00011011",	-- ...##.##
		1954 =>	"00011011",	-- ...##.##
		1955 =>	"00011000",	-- ...##...
		1956 =>	"00011000",	-- ...##...
		1957 =>	"00011000",	-- ...##...
		1958 =>	"00011000",	-- ...##...
		1959 =>	"00011000",	-- ...##...

		-- char 0xf5='\xf5
		1960 =>	"00011000",	-- ...##...
		1961 =>	"00011000",	-- ...##...
		1962 =>	"00011000",	-- ...##...
		1963 =>	"00011000",	-- ...##...
		1964 =>	"00011000",	-- ...##...
		1965 =>	"11011000",	-- ##.##...
		1966 =>	"11011000",	-- ##.##...
		1967 =>	"01110000",	-- .###....

		-- char 0xf6='\xf6
		1968 =>	"00110000",	-- ..##....
		1969 =>	"00110000",	-- ..##....
		1970 =>	"00000000",	-- ........
		1971 =>	"11111100",	-- ######..
		1972 =>	"00000000",	-- ........
		1973 =>	"00110000",	-- ..##....
		1974 =>	"00110000",	-- ..##....
		1975 =>	"00000000",	-- ........

		-- char 0xf7='\xf7
		1976 =>	"00000000",	-- ........
		1977 =>	"01110110",	-- .###.##.
		1978 =>	"11011100",	-- ##.###..
		1979 =>	"00000000",	-- ........
		1980 =>	"01110110",	-- .###.##.
		1981 =>	"11011100",	-- ##.###..
		1982 =>	"00000000",	-- ........
		1983 =>	"00000000",	-- ........

		-- char 0xf8='\xf8
		1984 =>	"00111000",	-- ..###...
		1985 =>	"01101100",	-- .##.##..
		1986 =>	"01101100",	-- .##.##..
		1987 =>	"00111000",	-- ..###...
		1988 =>	"00000000",	-- ........
		1989 =>	"00000000",	-- ........
		1990 =>	"00000000",	-- ........
		1991 =>	"00000000",	-- ........

		-- char 0xf9='\xf9
		1992 =>	"00000000",	-- ........
		1993 =>	"00000000",	-- ........
		1994 =>	"00000000",	-- ........
		1995 =>	"00011000",	-- ...##...
		1996 =>	"00011000",	-- ...##...
		1997 =>	"00000000",	-- ........
		1998 =>	"00000000",	-- ........
		1999 =>	"00000000",	-- ........

		-- char 0xfa='\xfa
		2000 =>	"00000000",	-- ........
		2001 =>	"00000000",	-- ........
		2002 =>	"00000000",	-- ........
		2003 =>	"00000000",	-- ........
		2004 =>	"00011000",	-- ...##...
		2005 =>	"00000000",	-- ........
		2006 =>	"00000000",	-- ........
		2007 =>	"00000000",	-- ........

		-- char 0xfb='\xfb
		2008 =>	"00001111",	-- ....####
		2009 =>	"00001100",	-- ....##..
		2010 =>	"00001100",	-- ....##..
		2011 =>	"00001100",	-- ....##..
		2012 =>	"11101100",	-- ###.##..
		2013 =>	"01101100",	-- .##.##..
		2014 =>	"00111100",	-- ..####..
		2015 =>	"00011100",	-- ...###..

		-- char 0xfc='\xfc
		2016 =>	"01111000",	-- .####...
		2017 =>	"01101100",	-- .##.##..
		2018 =>	"01101100",	-- .##.##..
		2019 =>	"01101100",	-- .##.##..
		2020 =>	"01101100",	-- .##.##..
		2021 =>	"00000000",	-- ........
		2022 =>	"00000000",	-- ........
		2023 =>	"00000000",	-- ........

		-- char 0xfd='\xfd
		2024 =>	"01110000",	-- .###....
		2025 =>	"00011000",	-- ...##...
		2026 =>	"00110000",	-- ..##....
		2027 =>	"01100000",	-- .##.....
		2028 =>	"01111000",	-- .####...
		2029 =>	"00000000",	-- ........
		2030 =>	"00000000",	-- ........
		2031 =>	"00000000",	-- ........

		-- char 0xfe='\xfe
		2032 =>	"00000000",	-- ........
		2033 =>	"00000000",	-- ........
		2034 =>	"00111100",	-- ..####..
		2035 =>	"00111100",	-- ..####..
		2036 =>	"00111100",	-- ..####..
		2037 =>	"00111100",	-- ..####..
		2038 =>	"00000000",	-- ........
		2039 =>	"00000000",	-- ........

		-- char 0xff='\xff
		2040 =>	"00000000",	-- ........
		2041 =>	"00000000",	-- ........
		2042 =>	"00000000",	-- ........
		2043 =>	"00000000",	-- ........
		2044 =>	"00000000",	-- ........
		2045 =>	"00000000",	-- ........
		2046 =>	"00000000",	-- ........
		2047 =>	"00000000",	-- ........
	others => (others => '0')
    );

end font8x8_xark;
