-- dual_config.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity dual_config is
	port (
		avmm_rcv_address   : in  std_logic_vector(2 downto 0)  := (others => '0'); -- avalon.address
		avmm_rcv_read      : in  std_logic                     := '0';             --       .read
		avmm_rcv_writedata : in  std_logic_vector(31 downto 0) := (others => '0'); --       .writedata
		avmm_rcv_write     : in  std_logic                     := '0';             --       .write
		avmm_rcv_readdata  : out std_logic_vector(31 downto 0);                    --       .readdata
		clk                : in  std_logic                     := '0';             --    clk.clk
		nreset             : in  std_logic                     := '0'              -- nreset.reset_n
	);
end entity dual_config;

architecture rtl of dual_config is
	component altera_dual_boot is
		generic (
			INTENDED_DEVICE_FAMILY : string  := "";
			CONFIG_CYCLE           : integer := 28;
			RESET_TIMER_CYCLE      : integer := 40
		);
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			nreset             : in  std_logic                     := 'X';             -- reset_n
			avmm_rcv_address   : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avmm_rcv_read      : in  std_logic                     := 'X';             -- read
			avmm_rcv_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avmm_rcv_write     : in  std_logic                     := 'X';             -- write
			avmm_rcv_readdata  : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component altera_dual_boot;

begin

	dual_boot_0 : component altera_dual_boot
		generic map (
			INTENDED_DEVICE_FAMILY => "MAX 10",
			CONFIG_CYCLE           => 9,
			RESET_TIMER_CYCLE      => 13
		)
		port map (
			clk                => clk,                --    clk.clk
			nreset             => nreset,             -- nreset.reset_n
			avmm_rcv_address   => avmm_rcv_address,   -- avalon.address
			avmm_rcv_read      => avmm_rcv_read,      --       .read
			avmm_rcv_writedata => avmm_rcv_writedata, --       .writedata
			avmm_rcv_write     => avmm_rcv_write,     --       .write
			avmm_rcv_readdata  => avmm_rcv_readdata   --       .readdata
		);

end architecture rtl; -- of dual_config
