library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package bootloader is
  type boot_block_type is array(0 to 511) of std_logic_vector(7 downto 0);

constant boot_block : boot_block_type := (
	x"13", x"07", x"07", x"ff", x"23", x"26", x"17", x"00", 
	x"23", x"24", x"27", x"00", x"23", x"22", x"37", x"00", 
	x"13", x"00", x"00", x"00", x"13", x"0b", x"00", x"00", 
	x"13", x"0a", x"00", x"00", x"37", x"1f", x"72", x"76", 
	x"b7", x"3e", x"3e", x"20", x"37", x"0e", x"00", x"08", 
	x"93", x"0b", x"30", x"00", x"93", x"0d", x"00", x"06", 
	x"13", x"0d", x"50", x"00", x"93", x"0c", x"00", x"04", 
	x"13", x"0c", x"f0", x"01", x"13", x"09", x"00", x"00", 
	x"93", x"08", x"df", x"a0", x"83", x"00", x"10", x"f2", 
	x"93", x"f9", x"40", x"00", x"e3", x"9c", x"09", x"fe", 
	x"23", x"00", x"10", x"f3", x"93", x"d8", x"88", x"40", 
	x"e3", x"96", x"08", x"fe", x"63", x"1a", x"09", x"02", 
	x"13", x"09", x"f0", x"ff", x"93", x"88", x"3e", x"23", 
	x"6f", x"f0", x"df", x"fd", x"13", x"08", x"00", x"00", 
	x"93", x"08", x"00", x"00", x"6f", x"00", x"80", x"06", 
	x"93", x"09", x"f0", x"0f", x"93", x"08", x"f0", x"ff", 
	x"93", x"0a", x"20", x"00", x"6f", x"00", x"00", x"02", 
	x"13", x"0b", x"08", x"00", x"6f", x"00", x"80", x"12", 
	x"93", x"09", x"f0", x"0f", x"93", x"08", x"f0", x"ff", 
	x"93", x"0a", x"20", x"00", x"93", x"00", x"20", x"00", 
	x"63", x"de", x"08", x"02", x"73", x"28", x"10", x"c0", 
	x"33", x"79", x"c8", x"01", x"63", x"06", x"09", x"00", 
	x"13", x"09", x"f0", x"0f", x"6f", x"00", x"80", x"00", 
	x"13", x"09", x"00", x"00", x"13", x"51", x"38", x"41", 
	x"93", x"71", x"f8", x"0f", x"13", x"71", x"f1", x"0f", 
	x"63", x"56", x"31", x"00", x"13", x"49", x"f9", x"00", 
	x"6f", x"00", x"00", x"01", x"13", x"49", x"09", x"0f", 
	x"6f", x"00", x"80", x"00", x"13", x"59", x"8a", x"40", 
	x"a3", x"08", x"20", x"f1", x"83", x"01", x"10", x"f2", 
	x"13", x"f9", x"11", x"00", x"e3", x"0a", x"09", x"fa", 
	x"03", x"09", x"00", x"f2", x"63", x"d6", x"08", x"02", 
	x"13", x"01", x"d9", x"fa", x"e3", x"08", x"01", x"f6", 
	x"93", x"01", x"39", x"ff", x"e3", x"8c", x"01", x"f2", 
	x"63", x"58", x"2c", x"07", x"03", x"08", x"10", x"f2", 
	x"13", x"78", x"48", x"00", x"e3", x"1c", x"08", x"fe", 
	x"23", x"00", x"20", x"f3", x"6f", x"f0", x"5f", x"f8", 
	x"13", x"01", x"69", x"ff", x"e3", x"fa", x"2b", x"f4", 
	x"13", x"18", x"48", x"00", x"63", x"d6", x"2d", x"01", 
	x"13", x"09", x"09", x"fe", x"6f", x"00", x"80", x"00", 
	x"63", x"d6", x"2c", x"01", x"13", x"09", x"99", x"fc", 
	x"6f", x"00", x"80", x"00", x"13", x"09", x"09", x"fd", 
	x"93", x"88", x"18", x"00", x"33", x"68", x"09", x"01", 
	x"13", x"89", x"f8", x"ff", x"63", x"1e", x"09", x"02", 
	x"93", x"01", x"98", x"ff", x"63", x"e2", x"30", x"02", 
	x"37", x"01", x"00", x"08", x"b7", x"01", x"01", x"00", 
	x"33", x"77", x"2b", x"00", x"33", x"67", x"37", x"00", 
	x"93", x"00", x"00", x"00", x"67", x"00", x"0b", x"00", 
	x"13", x"08", x"00", x"00", x"6f", x"f0", x"5f", x"f2", 
	x"e3", x"cc", x"0b", x"ff", x"93", x"19", x"18", x"00", 
	x"93", x"89", x"59", x"00", x"6f", x"f0", x"df", x"fe", 
	x"13", x"81", x"d8", x"ff", x"63", x"18", x"01", x"00", 
	x"13", x"18", x"18", x"00", x"b3", x"8a", x"0a", x"01", 
	x"6f", x"f0", x"9f", x"fd", x"e3", x"5e", x"3d", x"ef", 
	x"63", x"9a", x"38", x"01", x"13", x"0a", x"08", x"00", 
	x"e3", x"0c", x"0b", x"ec", x"93", x"89", x"08", x"00", 
	x"6f", x"f0", x"9f", x"ee", x"e3", x"d2", x"19", x"ef", 
	x"13", x"f9", x"18", x"00", x"e3", x"0e", x"09", x"ec", 
	x"e3", x"dc", x"58", x"ed", x"23", x"00", x"0a", x"01", 
	x"13", x"0a", x"1a", x"00", x"6f", x"f0", x"df", x"ec", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	others => (others => '0')
    );

end bootloader;
