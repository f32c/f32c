library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package bootloader is
  type boot_block_type is array(0 to 511) of std_logic_vector(7 downto 0);

constant boot_block : boot_block_type := (
	x"13", x"01", x"01", x"fe", x"23", x"2e", x"11", x"00", 
	x"23", x"2c", x"81", x"00", x"23", x"2a", x"91", x"00", 
	x"23", x"28", x"21", x"01", x"23", x"26", x"31", x"01", 
	x"23", x"24", x"41", x"01", x"23", x"22", x"51", x"01", 
	x"13", x"00", x"00", x"00", x"13", x"08", x"00", x"00", 
	x"93", x"05", x"00", x"00", x"93", x"07", x"00", x"00", 
	x"37", x"13", x"72", x"76", x"b7", x"33", x"3e", x"20", 
	x"37", x"0e", x"00", x"08", x"93", x"08", x"30", x"00", 
	x"93", x"0e", x"00", x"06", x"13", x"0f", x"10", x"00", 
	x"93", x"0f", x"50", x"00", x"93", x"00", x"00", x"04", 
	x"13", x"04", x"30", x"05", x"93", x"04", x"d0", x"00", 
	x"13", x"09", x"f0", x"01", x"13", x"0a", x"00", x"00", 
	x"13", x"07", x"d3", x"a0", x"03", x"06", x"10", x"f2", 
	x"93", x"12", x"d6", x"01", x"e3", x"cc", x"02", x"fe", 
	x"23", x"00", x"e0", x"f2", x"13", x"57", x"87", x"40", 
	x"33", x"65", x"47", x"01", x"63", x"18", x"05", x"00", 
	x"13", x"0a", x"f0", x"ff", x"13", x"87", x"33", x"23", 
	x"6f", x"f0", x"df", x"fd", x"e3", x"1c", x"07", x"fc", 
	x"13", x"05", x"20", x"00", x"13", x"06", x"f0", x"0f", 
	x"13", x"07", x"f0", x"ff", x"93", x"09", x"05", x"00", 
	x"13", x"da", x"85", x"40", x"63", x"5e", x"07", x"02", 
	x"f3", x"27", x"10", x"c0", x"b3", x"f6", x"c7", x"01", 
	x"b3", x"3a", x"d0", x"00", x"b3", x"02", x"50", x"41", 
	x"93", x"f6", x"f2", x"0f", x"93", x"d2", x"37", x"41", 
	x"93", x"fa", x"f7", x"0f", x"93", x"f2", x"f2", x"0f", 
	x"63", x"d6", x"52", x"01", x"93", x"c6", x"f6", x"00", 
	x"6f", x"00", x"80", x"00", x"93", x"c6", x"06", x"0f", 
	x"a3", x"08", x"d0", x"f0", x"6f", x"00", x"80", x"00", 
	x"a3", x"08", x"40", x"f1", x"83", x"0a", x"10", x"f2", 
	x"93", x"92", x"fa", x"01", x"e3", x"dc", x"02", x"fa", 
	x"03", x"0a", x"00", x"f2", x"63", x"5c", x"07", x"02", 
	x"63", x"18", x"8a", x"00", x"93", x"07", x"00", x"00", 
	x"13", x"07", x"00", x"00", x"6f", x"f0", x"df", x"f9", 
	x"e3", x"0a", x"9a", x"f4", x"93", x"07", x"00", x"00", 
	x"e3", x"58", x"49", x"f9", x"83", x"07", x"10", x"f2", 
	x"93", x"96", x"d7", x"01", x"e3", x"cc", x"06", x"fe", 
	x"23", x"00", x"40", x"f3", x"93", x"07", x"00", x"00", 
	x"6f", x"f0", x"9f", x"f7", x"93", x"06", x"6a", x"ff", 
	x"e3", x"f0", x"d8", x"f6", x"93", x"9a", x"47", x"00", 
	x"63", x"d6", x"4e", x"01", x"13", x"0a", x"0a", x"fe", 
	x"6f", x"00", x"00", x"01", x"93", x"07", x"0a", x"fd", 
	x"b3", x"e7", x"57", x"01", x"63", x"d6", x"40", x"01", 
	x"93", x"02", x"9a", x"fc", x"b3", x"e7", x"52", x"01", 
	x"13", x"07", x"17", x"00", x"63", x"1c", x"e7", x"03", 
	x"93", x"8a", x"97", x"ff", x"63", x"e0", x"59", x"03", 
	x"37", x"04", x"00", x"08", x"b7", x"04", x"01", x"00", 
	x"33", x"71", x"88", x"00", x"33", x"61", x"91", x"00", 
	x"93", x"00", x"00", x"00", x"67", x"00", x"08", x"00", 
	x"6f", x"f0", x"5f", x"fa", x"e3", x"c0", x"f8", x"fa", 
	x"93", x"92", x"17", x"00", x"13", x"86", x"52", x"00", 
	x"6f", x"f0", x"5f", x"f9", x"63", x"18", x"17", x"01", 
	x"93", x"96", x"17", x"00", x"33", x"05", x"d5", x"00", 
	x"6f", x"f0", x"5f", x"f8", x"e3", x"de", x"cf", x"ee", 
	x"63", x"1c", x"c7", x"00", x"93", x"85", x"07", x"00", 
	x"13", x"06", x"07", x"00", x"e3", x"16", x"08", x"ee", 
	x"13", x"88", x"07", x"00", x"6f", x"f0", x"5f", x"ee", 
	x"e3", x"50", x"e6", x"ee", x"13", x"1a", x"f7", x"01", 
	x"e3", x"5c", x"0a", x"ec", x"e3", x"5a", x"a7", x"ec", 
	x"23", x"80", x"f5", x"00", x"93", x"85", x"15", x"00", 
	x"6f", x"f0", x"9f", x"ec", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00", 
	others => (others => '0')
    );

end bootloader;
