library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

package bootloader is
  type boot_block_type is array(0 to 127) of std_logic_vector(7 downto 0);

constant boot_0 : boot_block_type := ( -- LSB bytes of 32-bit words
	x"00", x"21", x"21", x"66", x"3e", x"00", x"01", x"03", 
	x"53", x"0d", x"21", x"0d", x"21", x"04", x"fd", x"00", 
	x"20", x"03", x"25", x"04", x"00", x"ff", x"0c", x"32", 
	x"f3", x"ff", x"ff", x"02", x"1b", x"00", x"00", x"24", 
	x"02", x"21", x"ff", x"c3", x"ff", x"ff", x"2a", x"03", 
	x"00", x"2c", x"0f", x"f0", x"11", x"21", x"01", x"ec", 
	x"00", x"20", x"11", x"f6", x"05", x"00", x"21", x"21", 
	x"2c", x"03", x"cf", x"20", x"df", x"21", x"21", x"04", 
	x"fd", x"00", x"1c", x"20", x"04", x"05", x"00", x"ff", 
	x"ff", x"1e", x"02", x"61", x"03", x"d0", x"53", x"e0", 
	x"41", x"03", x"25", x"c9", x"25", x"01", x"11", x"f9", 
	x"03", x"09", x"04", x"00", x"10", x"24", x"21", x"08", 
	x"25", x"1c", x"21", x"fd", x"00", x"21", x"61", x"05", 
	x"04", x"06", x"21", x"61", x"21", x"ae", x"00", x"06", 
	x"2a", x"02", x"21", x"21", x"1c", x"21", x"a5", x"01", 
	x"a3", x"2a", x"a1", x"00", x"00", x"1c", x"01", x"00",
	others => (others => '0')
);

constant boot_1 : boot_block_type := (
	x"00", x"40", x"30", x"33", x"20", x"08", x"00", x"00", 
	x"00", x"00", x"c8", x"0a", x"ff", x"00", x"ff", x"00", 
	x"ff", x"1a", x"48", x"00", x"00", x"ff", x"00", x"63", 
	x"ff", x"00", x"ff", x"00", x"00", x"00", x"48", x"c8", 
	x"00", x"20", x"00", x"cc", x"00", x"00", x"48", x"00", 
	x"00", x"00", x"00", x"00", x"ff", x"ff", x"00", x"ff", 
	x"00", x"ff", x"00", x"ff", x"00", x"00", x"10", x"18", 
	x"00", x"22", x"ff", x"00", x"ff", x"10", x"ff", x"00", 
	x"ff", x"00", x"00", x"ff", x"00", x"00", x"49", x"00", 
	x"ff", x"00", x"00", x"00", x"00", x"ff", x"00", x"ff", 
	x"00", x"00", x"10", x"ff", x"10", x"00", x"00", x"ff", 
	x"00", x"00", x"00", x"80", x"00", x"e8", x"f8", x"00", 
	x"e8", x"00", x"10", x"ff", x"00", x"28", x"00", x"00", 
	x"00", x"00", x"10", x"00", x"38", x"ff", x"00", x"00", 
	x"c8", x"00", x"30", x"40", x"00", x"28", x"ff", x"00", 
	x"ff", x"48", x"ff", x"00", x"00", x"00", x"00", x"00",
	others => (others => '0')
);

constant boot_2 : boot_block_type := (
	x"00", x"00", x"00", x"0a", x"0b", x"0c", x"0d", x"0e", 
	x"0f", x"18", x"00", x"43", x"05", x"a7", x"e0", x"00", 
	x"03", x"03", x"79", x"20", x"00", x"19", x"00", x"63", 
	x"60", x"05", x"03", x"07", x"61", x"00", x"02", x"4c", 
	x"20", x"00", x"04", x"02", x"49", x"39", x"29", x"20", 
	x"00", x"00", x"84", x"84", x"04", x"04", x"99", x"20", 
	x"00", x"04", x"61", x"89", x"8f", x"00", x"00", x"00", 
	x"00", x"06", x"98", x"99", x"20", x"00", x"02", x"42", 
	x"40", x"00", x"00", x"04", x"39", x"20", x"02", x"05", 
	x"03", x"00", x"07", x"82", x"40", x"82", x"00", x"84", 
	x"99", x"20", x"49", x"84", x"89", x"63", x"6d", x"59", 
	x"24", x"80", x"49", x"04", x"05", x"04", x"00", x"00", 
	x"a5", x"00", x"00", x"20", x"00", x"42", x"00", x"a5", 
	x"6e", x"a9", x"42", x"00", x"e2", x"20", x"00", x"65", 
	x"a3", x"00", x"40", x"40", x"00", x"60", x"20", x"64", 
	x"80", x"67", x"20", x"00", x"c2", x"00", x"c6", x"00",
	others => (others => '0')
);

constant boot_3 : boot_block_type := ( -- MSB bytes of 32-bit words
	x"00", x"00", x"00", x"3c", x"3c", x"3c", x"24", x"24", 
	x"24", x"24", x"00", x"25", x"80", x"30", x"14", x"00", 
	x"a0", x"00", x"00", x"15", x"00", x"24", x"08", x"25", 
	x"14", x"24", x"24", x"24", x"04", x"00", x"40", x"00", 
	x"13", x"00", x"24", x"00", x"30", x"33", x"03", x"11", 
	x"00", x"08", x"38", x"38", x"a0", x"80", x"30", x"13", 
	x"00", x"80", x"04", x"24", x"14", x"00", x"00", x"00", 
	x"08", x"00", x"10", x"28", x"17", x"00", x"80", x"30", 
	x"14", x"00", x"08", x"a0", x"2d", x"13", x"00", x"24", 
	x"24", x"08", x"24", x"28", x"14", x"24", x"08", x"24", 
	x"28", x"17", x"00", x"24", x"00", x"24", x"14", x"24", 
	x"2f", x"10", x"28", x"3c", x"3c", x"01", x"00", x"01", 
	x"03", x"08", x"00", x"11", x"00", x"00", x"08", x"24", 
	x"14", x"28", x"00", x"08", x"00", x"15", x"00", x"14", 
	x"00", x"15", x"00", x"00", x"08", x"00", x"13", x"30", 
	x"10", x"00", x"11", x"00", x"a0", x"08", x"24", x"00",
	others => (others => '0')
);

end bootloader;
