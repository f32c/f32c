--
-- Copyright 2008, 2010 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
--

-- $Id$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Xilinx libraries
library UNISIM;
use UNISIM.VComponents.all;

entity bram is
	generic(
		mem_type: string := "big"
	);
	port(
		clk: in std_logic;
		imem_addr: in std_logic_vector(31 downto 2);
		imem_data_out: out std_logic_vector(31 downto 0);
		imem_addr_strobe: in std_logic;
		imem_data_ready: out std_logic;
		dmem_addr: in std_logic_vector(31 downto 2);
		dmem_data_in: in std_logic_vector(31 downto 0);
		dmem_data_out: out std_logic_vector(31 downto 0);
		dmem_byte_we: in std_logic_vector(3 downto 0);
		dmem_addr_strobe: in std_logic;
		dmem_data_ready: out std_logic
	);
end bram;

architecture Behavioral of bram is
	signal dmem_wait_cycle, dmem_must_wait, dmem_we: std_logic;
	signal dmem_data_read, dmem_write_out: std_logic_vector(31 downto 0);
	signal dmem_bram_cs: std_logic;
begin
	
	imem_data_ready <= '1';
	dmem_data_out <= dmem_data_read; -- shut up compiler errors
	
	-- 32-bit wide memory with wait state insertion on byte / half word writes
	small_mem:
	if mem_type = "small" generate
	begin
	
	dmem_data_ready <= not dmem_must_wait;
	
	-- We need a read followed by a write cycle if storing a byte or half a word, so
	-- insert a wait state in such cases
	dmem_must_wait <= '1' when dmem_wait_cycle = '0' and dmem_byte_we /= "0000" and
		dmem_byte_we /= "1111" and dmem_addr_strobe = '1' else '0';
	
	process(clk, dmem_must_wait)
	begin
		if rising_edge(clk) then
			if dmem_wait_cycle = '0' and dmem_must_wait = '1' then
				dmem_wait_cycle <= '1';
			else
				dmem_wait_cycle <= '0';
			end if;
		end if;
	end process;
	
	dmem_we <= '1' when dmem_byte_we /= "0000" and dmem_must_wait = '0' else '0';
	dmem_write_out(7 downto 0) <= dmem_data_in(7 downto 0) when
		dmem_byte_we(0) = '1' else dmem_data_read(7 downto 0);
	dmem_write_out(15 downto 8) <= dmem_data_in(15 downto 8) when
		dmem_byte_we(1) = '1' else dmem_data_read(15 downto 8);
	dmem_write_out(23 downto 16) <= dmem_data_in(23 downto 16) when
		dmem_byte_we(2) = '1' else dmem_data_read(23 downto 16);
	dmem_write_out(31 downto 24) <= dmem_data_in(31 downto 24) when
		dmem_byte_we(3) = '1' else dmem_data_read(31 downto 24);
	
	dmem_bram_cs <= dmem_addr_strobe;
	dmem: RAMB16_S36_S36
		generic map(
			INIT_00 => x"000000001000fff98f7a00043c1be0000c0002fc3c1d0001379c8d803c1c0000",
			INIT_01 => x"000b508224cbfffc144000153042000300a41025008038211440001728c20004",
			INIT_02 => x"1509fffb2508000400a818218c44000000e81021000040210002488025420001",
			INIT_03 => x"00a2282101633023000a188000021080244200010002108224c2fffcac640000",
			INIT_04 => x"1cc0fffba0a2000024e7000124c6ffff90e200000000000018c0000700e23821",
			INIT_05 => x"1440001730820003008038211440001828c200040000000003e0000824a50001",
			INIT_06 => x"00021c00000420802524000100451021000a48820005120024cafffc00051600",
			INIT_07 => x"0002108224c2fffc1488fffd24840004ac83000000e020210062182100e44021",
			INIT_08 => x"000216030005160018c0000600e2382101433023000210800009188024420001",
			INIT_09 => x"1040000a308200030000000003e0000824e700011cc0fffda0e2000024c6ffff",
			INIT_0A => x"246300011440fffd808200002484000100001821104000058082000000002821",
			INIT_0B => x"248400048c85000000052a031440000330620003000018210060102103e00008",
			INIT_0C => x"00001821108000080060102103e000082463ffff246300011440fff930a200ff",
			INIT_0D => x"03e00008000000001480fffa0004204000641821000528421040000230a20001",
			INIT_0E => x"012a2825240b00200800007a0000182100052fc00000402100a0382100601021",
			INIT_0F => x"1440fff724630001000550420085102b00024f8030e2000200073842106b0011",
			INIT_10 => x"012a28253508000100852023000000001040fff32ce2000210a0fff500084040",
			INIT_11 => x"8f8480b00100102103e00008acc400000000000010c0000200073842146bfff1",
			INIT_12 => x"0c00007134a5f31d3c0500013444d9243c02075bafbf001c1480000327bdffe0",
			INIT_13 => x"00c33021000719c00007314000a3282300022980000218808fa7001027a60010",
			INIT_14 => x"0062182100031880008720210086202300651823000621000005188000a22823",
			INIT_15 => x"3442ffff3c027fff8fbf001c04610004004318230003188000441023000410c0",
			INIT_16 => x"afbf0024afb0001827bdffd827bd002003e00008af8380b00060102100621821",
			INIT_17 => x"00c0882127b20010080000c00200882100a0802104800024afb1001cafb20020",
			INIT_18 => x"00022e0024420030262600018fa2001000402021024030210c0000712405000a",
			INIT_19 => x"02201821080000d18fbf00241040000c0211102ba22500001480fff500052e03",
			INIT_1A => x"1440fff80203102b2463ffffa062000026100001a20500008202000080650000",
			INIT_1B => x"2402002d27bd002803e000088fb000188fb1001c8fb2002000c010218fbf0024",
			INIT_1C => x"24080008080000ec0000182124a5000124b00001080000bc00042023a0a20000",
			INIT_1D => x"2842000a24460030244700570004170224a500011068000ba0a7ffff24630001",
			INIT_1E => x"0000000003e0000824a500011468fff7a0a6ffff24630001000421001040fff7",
			INIT_1F => x"3403c350000088211080000b00802821afb00014afbf001cafb1001827bdffe0",
			INIT_20 => x"3062000114a0fffb000528400085202100031842104000023062000100002021",
			INIT_21 => x"0043102400821026af8480b88f8380108f8280b48f6400008f70000400808821",
			INIT_22 => x"8f620004000000000c000128af8480b48fbf001c1460000d0064182410400004",
			INIT_23 => x"27bd002003e000088fb000148fb100188fbf001c1440ffef0051102a00501023",
			INIT_24 => x"00000000000000000000000027bd002003e000088fb000148fb1001824020001",
			INIT_25 => x"00002821344420003c02004eafb000001440002fafb1000427bdfff88f8280a0",
			INIT_26 => x"8f6200048f630004af67000caf66000824090003000040212407000224060038",
			INIT_27 => x"004310238f6200048f630004af68000c000000001440fffc0044102a00431023",
			INIT_28 => x"24030002af6200082402000c14a9ffef24a50001000000001440fffc0044102a",
			INIT_29 => x"1440fffc0044102a004310238f620004344488003c0200138f630004af63000c",
			INIT_2A => x"0044102a004310238f620004344488003c0200138f630004af62000c00000000",
			INIT_2B => x"304a0001000210c38f8780b48f8980148f620000af8280a0240200011440fffc",
			INIT_2C => x"2418f9ff2411020024100400240f0600240e0003240d00010000c821278b80c0",
			INIT_2D => x"240300941322000424020002144000582b220002240300c0132d0009240c0004",
			INIT_2E => x"8f6200048f630004af62000c24020002af63000800001821240300d4132e0002",
			INIT_2F => x"004310238f6200048f630004af62000c000000001440fffc2842138800431023",
			INIT_30 => x"000000001040002a010b102b256b001401604021000000001440fffc28421388",
			INIT_31 => x"1440000528620061000632031140000800031e0300061e00000028218d060000",
			INIT_32 => x"108f0022304406008f62000000031e0300021e002462ffe0104000032862007b",
			INIT_33 => x"004310238f6200048f630004af6e000caf6300080082382500f8102430e20600",
			INIT_34 => x"28421388004310238f6200048f630004af6d000c000000001440fffc28421388",
			INIT_35 => x"1440ffd8010b102b250800040000000014acffde24a50001000000001440fffc",
			INIT_36 => x"af8780b4af8980148fb000008fb1000400000000172cffb62739000100000000",
			INIT_37 => x"2c4200012922ffc100f810241451ffdd000000001050000727bd000803e00008",
			INIT_38 => x"08000173240300801320ffad01224821080001992922003f0122482308000199",
			INIT_39 => x"afb50024afbf002cafb6002827bdffd000000000000000000000000000001821",
			INIT_3A => x"00a0b0211080003300803021afb00010afb10014afb20018afb3001cafb40020",
			INIT_3B => x"004410210006108000062100af620000af8280a400a21025304200f08f8280a4",
			INIT_3C => x"000210838f620000240600140c00002b24050020028020210043a021278380e8",
			INIT_3D => x"2415001500008821006490212784806c00621823000210c00002194030420001",
			INIT_3E => x"8fbf002c265200081635fffa263100071440000d02c21024029198218e420000",
			INIT_3F => x"03e000088fb000108fb100148fb200188fb3001c8fb400208fb500248fb60028"
		)
		port map(
			DIA => dmem_write_out, DIB => x"ffffffff",
			DOA => dmem_data_read, DOB => imem_data_out,
			ADDRA => dmem_addr(10 downto 2),	ADDRB => imem_addr(10 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_we, WEB => '0', DIPA => x"f", DIPB => x"f"
		);

	end generate; -- small_mem
	
	big_mem:
	if mem_type /= "small" generate
	begin
	
	dmem_data_ready <= '1';
	dmem_write_out <= dmem_data_in;
	dmem_bram_cs <= dmem_addr_strobe;
		
	dmem_0: RAMB16_S9_S9
		generic map(
			INIT_00 => x"212380800182fc00fb0421002121800182fc15032521170400f90400fc018000",
			INIT_01 => x"82fcfd0400212121008001218200fc001703211804000801fb0001ff00000721",
			INIT_02 => x"040003030321210801fd0001210500210a03000801fd00ff0300062123808001",
			INIT_03 => x"f701422b8002421125207a21c02121210800fa402142020121082108ff01f9ff",
			INIT_04 => x"21c0402380801010711d01245b1c03e0b0210800000242f125012300f302f540",
			INIT_05 => x"2110c02121241c202418d82008b02121ffff1c04238023c02180212323008023",
			INIT_06 => x"2d2808181c202124f82bff000100000021d1240c2b00f503003001102121710a",
			INIT_07 => x"50210b21141c18e0000801f7ff0100f70a305702010bff0108ec210101bc2300",
			INIT_08 => x"200814181cef2a23040028b41c0d24042426b810b400042101fb402142020121",
			INIT_09 => x"2304040c00fc2a2304040c080321023821004e002f04f8a00000002008141801",
			INIT_0A => x"01c3b41400a001fc2a23040013040c00fc2a23040013040c02080cef0100fc2a",
			INIT_0B => x"2304040c00fc882304040c020821d4029404025802c00904ff000000030121c0",
			INIT_0C => x"2304040c082524002200000300e0037b0561030803002100002a2b142100fc88",
			INIT_0D => x"01c124dd00070808b414000400b60100d82b0400de0100fc882304040c00fc88",
			INIT_0E => x"21800000a425f0a42133211014181c20242c28d0000000217380ad21993f2399",
			INIT_0F => x"081014181c2024282c08fa070d2421001521216c23c040018300142b202121e8",
			INIT_10 => x"c04e1c2024282c212118001421d01880a4dc250f00a400f521082121214e0430",
			INIT_11 => x"07002138142c14fc2b1420142b20e8142b20d4a84d04b903a702920121082121",
			INIT_12 => x"23b526c32303000021213021082121284323214e002108212121144323214ec0",
			INIT_13 => x"a8ccac0121010830f814181c2024282c6400440024012171407d04030821a000",
			INIT_14 => x"40f802cca82ceedcf80ccca864700021300814181c2024282c000edcf808ccac",
			INIT_15 => x"f41421cc0121cc21b87004cca800f12cd8f4f8a8cc02ddf4f801cc21a80421e6",
			INIT_16 => x"14181c2024282c0ecc4001140ecc8321142370c01404cc0104cc212cc423f8c0",
			INIT_17 => x"1420c0e830f82314181c202428c0ff2c14a80ecc01a8a8cc210ec3008f30f864",
			INIT_18 => x"199cb4101418149c0605019c0d242610b4b8142bfc20142b20e8142b20d4142b",
			INIT_19 => x"6e70206f656c752000612075206f656e76206673736f2020000000b410181421",
			INIT_1A => x"6f7964206e7a6f206e636b6f447453725a6947006f4b655a6f696f5376566575",
			INIT_1B => x"02600458087d4c9a441f3cc934372800204010da08f4e0ccb8a43f0000006e67",
			INIT_1C => x"0000000000000000000000000000000000000000000000000380027804700868",
			INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(7 downto 0), DIB => x"ff",
			DOA => dmem_data_read(7 downto 0), DOB => imem_data_out(7 downto 0),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(0), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_1: RAMB16_S9_S9
		generic map(
			INIT_00 => x"283018100010ff00ff0018001040480050ff00001038000000ff00e002008d00",
			INIT_01 => x"10ffff00002018401c2000104812ff160000380000000000ff0000ff00000038",
			INIT_02 => x"00002a000018100000ff0000180000280000000000ff00ff1616003830101800",
			INIT_03 => x"ff0050104f003800280000182f4038100000ff201828000018001000ff00ff00",
			INIT_04 => x"301931282918000000f300d9070000ff80100000000038ff28002000ff00ff40",
			INIT_05 => x"88000088800000000000ff0000801018ff7f0000181810101818202018211828",
			INIT_06 => x"0000000000001000ff10ff0000000000180000001000ff2e2e00000020300000",
			INIT_07 => x"c3880028000000ff000000ffff0021ff000000170000ff000000180000002000",
			INIT_08 => x"0000000000ff10100000018000001800101080808000008800ff282018000020",
			INIT_09 => x"1000000000ff10100000000000400000282000000000ff800000000000000000",
			INIT_0A => x"00108080008000ff1010008800000000ff10100088000000000000ff0000ff10",
			INIT_0B => x"1000000000ff131000000000001800000000000000000000f90204060000c880",
			INIT_0C => x"10000000003810060006001e1eff0000000032001e1e2800000010004000ff13",
			INIT_0D => x"00ff10ff000000008080000000ff0000ff100000ff0000ff131000000000ff13",
			INIT_0E => x"1010210080100080b000300000000000000000ff000000180100ff4801004801",
			INIT_0F => x"00000000000000000000ff00001098000088908018101900100000000020a080",
			INIT_10 => x"80000000000000208800000010ff801880011000198000012800203020000000",
			INIT_11 => x"0000100000808080000000000000800000008080000000000000000028002030",
			INIT_12 => x"2000201720810000108880200028300080802000009000203028002828200088",
			INIT_13 => x"8001800020000000000000000000000000000000000030007801000000280c00",
			INIT_14 => x"1f0000018000ff05000001800002001000000000000000000000000500000180",
			INIT_15 => x"01802801002801200b0200018000ff00ff0100800100ff0100000128800080ff",
			INIT_16 => x"00000000000000000128008000012820802002208000010000012000ff200020",
			INIT_17 => x"000080ff00002000000000000020010080800001008080012000280000000000",
			INIT_18 => x"0380800280000080000000800010108080800000800000000080000000800000",
			INIT_19 => x"656c20726d6964500066736320726d6961506f656b6d416b0000008002000020",
			INIT_1A => x"776500206f65007a6f7200767500700061636f007661626164206e6c61750063",
			INIT_1B => x"000d000d00020d010d010d000d000d000dff0dfe0d0c0c0c0c0c000100000072",
			INIT_1C => x"000000000000000000000000000000000000000000000000000d000d000d000d",
			INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(15 downto 8), DIB => x"ff",
			DOA => dmem_data_read(15 downto 8), DOB => imem_data_out(15 downto 8),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(1), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_2: RAMB16_S9_S9
		generic map(
			INIT_00 => x"a2630a024202c2640908a844e80002420bcb4042a48040c200007a1b001d9c1c",
			INIT_01 => x"02c2888483e062e4020424450a05ca0540828040c200e0a5c0a2e7c6e200c0e2",
			INIT_02 => x"84850540620060e06340828400408200408200e0e7c0e2c60205c0e243020942",
			INIT_03 => x"4063058502e2076b2a0b00000500a060e0008004640540a2008060e0636340a2",
			INIT_04 => x"c30707a30202a7a600a5054402bf80bd8400e0c400c0076b2a08850040e2a008",
			INIT_05 => x"c0b20000a080b1b2bfb0bdbde08360624202bf614303440462038786650605a2",
			INIT_06 => x"02bde0b0b1b2c0bf40036362100502652000bf4011258005024226a240400005",
			INIT_07 => x"03008080b0bfb1bd00e0a568a663044042464704a568a763080000a5b00004a2",
			INIT_08 => x"bde0b0b1bf40515062000084bf606440438284838264708062a0058503406200",
			INIT_09 => x"43626368004044436263676609000706004402b040b1bd82000000bde0b0b102",
			INIT_0A => x"4a0287896282024044436244026362004044436244026363036202a9a5004044",
			INIT_0B => x"4362636200404243626362026300032e0322024022032d0c1811100f0e0d008b",
			INIT_0C => x"4362636e6382f8e28f44620302624062406206400306000600400b6b60004042",
			INIT_0D => x"4222f8510050bde08789b0b1002c3900400b0800aca50040424362636d004042",
			INIT_0E => x"4406066282a24282a08080b0b1b2b3b4b5bfb6bd000000000003202200222200",
			INIT_0F => x"e0b0b1b2b3b4b5b6bf52353140c2914215006484620202420262060005804383",
			INIT_10 => x"9500b2b3b4b5bf0080b150b043bd8204820062420582000060000040000050bd",
			INIT_11 => x"31535434109291840006050600058406000584822202220222022202a0000040",
			INIT_12 => x"82004404838544235451826000b04010100260005351006040a5a50502600011",
			INIT_13 => x"82008343404205bd00b0b1b2b3b4b5bf0462020040420000a505640600408404",
			INIT_14 => x"0400050084bf40040005008404006200bde0b0b1b2b3b4b5bf00400400050084",
			INIT_15 => x"108400000400000004000500840011bf40040084000540040010000084110040",
			INIT_16 => x"b0b1b2b3b4b5bfa500050485a50005008504000484050004050000bf40040004",
			INIT_17 => x"bf0584bdbd0044b0b1b2b3b4b50442bf8482a5000485820000a5020000bd0004",
			INIT_18 => x"0080850080bdbf84408284844043a28382850600840506000584060005840600",
			INIT_19 => x"20614e0061206a6f006f656e20006120726f726d6961756d0000008500bdbf00",
			INIT_1A => x"006c0072006c00750076006e62006c00640073006172006700427361726b0069",
			INIT_1B => x"0000000000000000000000000000000000ff00ff000000000000000000000065",
			INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(23 downto 16), DIB => x"ff",
			DOA => dmem_data_read(23 downto 16), DOB => imem_data_out(23 downto 16),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(2), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_3: RAMB16_S9_S9
		generic map(
			INIT_00 => x"00010000240024ac1525008c00000025002414300000142800108f3c0c3c373c",
			INIT_01 => x"00241424ac000000000025000000240014300014280003241ca0242490001800",
			INIT_02 => x"248c001430000003241480240010800010300003241ca0240000180001000024",
			INIT_03 => x"1424000000300010012408000000000003001400000010300010000324241430",
			INIT_04 => x"0000000000008f270c343c343caf14278f0103ac0010001401350000102c1000",
			INIT_05 => x"002708020004afafafaf272703af0000343c8f04000000000000000000000000",
			INIT_06 => x"2427038f8f8f008f140224a026a2828002088f1002a214000024268f00020c24",
			INIT_07 => x"34001000afafaf2700032414a0240010282424002410a02424080024240800a0",
			INIT_08 => x"27038f8f8f1400008f000caf8f1400100000af8f8f8f8f003014000000103000",
			INIT_09 => x"008f8faf001400008f8fafaf2400242400343caf14af278f00000027038f8f24",
			INIT_0A => x"30008f8f8faf241400008f343c8faf001400008f343c8faf24af241424001400",
			INIT_0B => x"008f8faf001428008f8faf24af002413241324142b2413242424242424240027",
			INIT_0C => x"008f8fafaf00003010308f0000241028142800110000008d0010012501001428",
			INIT_0D => x"2c29001400102703afaf8f8f00172700140125001424001428008f8faf001428",
			INIT_0E => x"000000afaf00308f001000afafafafafafafaf27000000000824130108290108",
			INIT_0F => x"038f8f8f8f8f8f8f8f2616261402028e2400002700000030008f240c24020027",
			INIT_10 => x"270cafafafafaf0200af8caf00272700af080030008f0008020c0200020c8e27",
			INIT_11 => x"328c023224278f270c2424240c2427240c24278f1624122412241224020c0200",
			INIT_12 => x"000c000000278c8e000027020c0200260002020c8e020c020002240002020c00",
			INIT_13 => x"af0caf2c002c2427088f8f8f8f8f8f8f24af24001030000c343c8f240c00243c",
			INIT_14 => x"240c240c8f8f14240c240c8f2408af0027038f8f8f8f8f8f8f0010240c240c8f",
			INIT_15 => x"248f000c24000c002408240c8f00168f14240c8f0c2414240c260c008f240014",
			INIT_16 => x"8f8f8f8f8f8f8f300c00248f300c00008f0208008f240c24240c008f14020c00",
			INIT_17 => x"af2427272708008f8f8f8f8f8f00308f8f8f300c248faf0c003000000c270824",
			INIT_18 => x"08afaf08af278faf1028248f1000008f8f8f240c2724240c2427240c2427240c",
			INIT_19 => x"6b7461006673656c00726d6952006673656b006120747400000000af08278f00",
			INIT_1A => x"006c006500650074006500697200690061007000636c007200726b76006f0063",
			INIT_1B => x"0000000000000000000000000000000000ff00ff000000000000000000000065",
			INIT_1C => x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1D => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(31 downto 24), DIB => x"ff",
			DOA => dmem_data_read(31 downto 24), DOB => imem_data_out(31 downto 24),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(3), WEB => '0', DIPA => "1", DIPB => "1"
		);
		
	end generate; -- big_mem
end Behavioral;
