--
-- Copyright 2008, 2010 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
--

-- $Id$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Xilinx libraries
library UNISIM;
use UNISIM.VComponents.all;

entity bram is
	generic(
		mem_type: string := "big"
	);
	port(
		clk: in std_logic;
		imem_addr: in std_logic_vector(31 downto 2);
		imem_data_out: out std_logic_vector(31 downto 0);
		imem_addr_strobe: in std_logic;
		imem_data_ready: out std_logic;
		dmem_addr: in std_logic_vector(31 downto 2);
		dmem_data_in: in std_logic_vector(31 downto 0);
		dmem_data_out: out std_logic_vector(31 downto 0);
		dmem_byte_we: in std_logic_vector(3 downto 0);
		dmem_addr_strobe: in std_logic;
		dmem_data_ready: out std_logic
	);
end bram;

architecture Behavioral of bram is
	signal dmem_wait_cycle, dmem_must_wait, dmem_we: std_logic;
	signal dmem_data_read, dmem_write_out: std_logic_vector(31 downto 0);
	signal dmem_bram_cs: std_logic;
begin
	
	imem_data_ready <= '1';
	dmem_data_out <= dmem_data_read; -- shut up compiler errors
	
	-- 32-bit wide memory with wait state insertion on byte / half word writes
	small_mem:
	if mem_type = "small" generate
	begin
	
	dmem_data_ready <= not dmem_must_wait;
	
	-- We need a read followed by a write cycle if storing a byte or half a word, so
	-- insert a wait state in such cases
	dmem_must_wait <= '1' when dmem_wait_cycle = '0' and dmem_byte_we /= "0000" and
		dmem_byte_we /= "1111" and dmem_addr_strobe = '1' else '0';
	
	process(clk, dmem_must_wait)
	begin
		if rising_edge(clk) then
			if dmem_wait_cycle = '0' and dmem_must_wait = '1' then
				dmem_wait_cycle <= '1';
			else
				dmem_wait_cycle <= '0';
			end if;
		end if;
	end process;
	
	dmem_we <= '1' when dmem_byte_we /= "0000" and dmem_must_wait = '0' else '0';
	dmem_write_out(7 downto 0) <= dmem_data_in(7 downto 0) when
		dmem_byte_we(0) = '1' else dmem_data_read(7 downto 0);
	dmem_write_out(15 downto 8) <= dmem_data_in(15 downto 8) when
		dmem_byte_we(1) = '1' else dmem_data_read(15 downto 8);
	dmem_write_out(23 downto 16) <= dmem_data_in(23 downto 16) when
		dmem_byte_we(2) = '1' else dmem_data_read(23 downto 16);
	dmem_write_out(31 downto 24) <= dmem_data_in(31 downto 24) when
		dmem_byte_we(3) = '1' else dmem_data_read(31 downto 24);
	
	dmem_bram_cs <= dmem_addr_strobe;
	dmem: RAMB16_S36_S36
		generic map(
			INIT_00 => x"00000000000000001000fffa3c1be0000c0002c03c1d0001379c8c903c1c0000",
			INIT_01 => x"24a500011cc0fffba0a200002484000124c6ffff908200000000000018c00007",
			INIT_02 => x"1cc0fffda085000024c6ffff00052e0300052e0018c000060000000003e00008",
			INIT_03 => x"80820000248400010000182110400005808200000000000003e0000824840001",
			INIT_04 => x"1040000230a2000100001821108000080060102103e00008246300011440fffd",
			INIT_05 => x"00a038210060102103e00008000000001480fffa000420400064182100052842",
			INIT_06 => x"00073842106b0011012a2825240b0020080000380000182100052fc000004021",
			INIT_07 => x"10a0fff5000840401440fff724630001000550420085102b00024f8030e20002",
			INIT_08 => x"00073842146bfff1012a28253508000100852023000000001040fff32ce20002",
			INIT_09 => x"1480000327bdffe08f8480ac0100102103e00008acc400000000000010c00002",
			INIT_0A => x"8fa7001027a600100c00002f34a5f31d3c0500013444d9243c02075bafbf001c",
			INIT_0B => x"0005188000a2282300c33021000719c00007314000a328230002298000021880",
			INIT_0C => x"00441023000410c0006218210003188000872021008620230065182300062100",
			INIT_0D => x"00601021006218213442ffff3c027fff8fbf001c046100040043182300031880",
			INIT_0E => x"afb1001cafb20020afbf0024afb0001827bdffd827bd002003e00008af8380ac",
			INIT_0F => x"0c00002f2405000a00c0882127b200100800007e0200882100a0802104800024",
			INIT_10 => x"1480fff500052e0300022e0024420030262600018fa200100040202102403021",
			INIT_11 => x"8202000080650000022018210800008f8fbf00241040000c0211102ba2250000",
			INIT_12 => x"00c010218fbf00241440fff80203102b2463ffffa062000026100001a2050000",
			INIT_13 => x"00042023a0a200002402002d27bd002803e000088fb000188fb1001c8fb20020",
			INIT_14 => x"a0a7ffff2463000124080008080000aa0000182124a5000124b000010800007a",
			INIT_15 => x"000421001040fff72842000a24460030244700570004170224a500011068000b",
			INIT_16 => x"afb1001827bdffe00000000003e0000824a500011468fff7a0a6ffff24630001",
			INIT_17 => x"30620001000020213403c350000088211080000b00802821afb00014afbf001c",
			INIT_18 => x"8f700004008088213062000114a0fffb00052840008520210003184210400002",
			INIT_19 => x"00641824104000040043102400821026af8480b88f8380108f8280b48f640000",
			INIT_1A => x"0051102a005010238f620004000000000c0000e4af8480b48fbf001c1460000d",
			INIT_1B => x"8fb100182402000127bd002003e000088fb000148fb100188fbf001c1440ffef",
			INIT_1C => x"afb20018afbf001c27bdffe08f8280980000000027bd002003e000088fb00014",
			INIT_1D => x"240700022406003800002821344420003c02004eafb000101440002fafb10014",
			INIT_1E => x"0044102a004310238f6200048f630004af67000caf6600082409000300004021",
			INIT_1F => x"1440fffc0044102a004310238f6200048f630004af68000c000000001440fffc",
			INIT_20 => x"8f630004af63000c24030002af6200082402000c14a9ffef24a5000100000000",
			INIT_21 => x"af62000c000000001440fffc0044102a004310238f620004344488003c020013",
			INIT_22 => x"240200011440fffc0044102a004310238f620004344488003c0200138f630004",
			INIT_23 => x"00042400278580de978280b88f8480b4278580d40c0000a28f640004af828098",
			INIT_24 => x"00004821304a0001000210c38f8780b48f8880b08f620000004420250c0000a2",
			INIT_25 => x"2419020024180400240d0600240c00032411000200008021240b0001279f80c0",
			INIT_26 => x"000000001440005129220002240200c0112b000924120004240f0014240ef9ff",
			INIT_27 => x"8f630004af71000caf62000800001021240200d4112c00022402009411310004",
			INIT_28 => x"8f6200048f630004af70000c000000001440fffc28421388004310238f620004",
			INIT_29 => x"0000282103e230210043102100091900000910801440fffc2842138800431023",
			INIT_2A => x"00021e002462ffe0104000032862007b144000052862006180c3000011400008",
			INIT_2B => x"af6300080044382500ee1024af8280b8108d0020304406008f62000000031e03",
			INIT_2C => x"af6b000c000000001440fffc28421388004310238f6200048f630004af6c000c",
			INIT_2D => x"14afffe024a50001000000001440fffc28421388004310238f6200048f630004",
			INIT_2E => x"8fb000108fb100148fb200188fbf001c000000001532ffc02529000124c60001",
			INIT_2F => x"1459ffde000000001058000730e2060027bd002003e00008af8780b4af8880b0",
			INIT_30 => x"010240210800015d2902003f010240230800015d2c4200012902ffc100ee1024",
			INIT_31 => x"afb50024afbf002cafb6002827bdffd0000010210800013d240200801120ffb4",
			INIT_32 => x"00a0b0211080003300803021afb00010afb10014afb20018afb3001cafb40020",
			INIT_33 => x"004410210006108000062100af620000af82809c00a21025304200f08f82809c",
			INIT_34 => x"000210838f620000240600140c00001224050020028020210043a021278380e8",
			INIT_35 => x"2415001500008821006490212784806800621823000210c00002194030420001",
			INIT_36 => x"8fbf002c265200081635fffa263100071440000d02c21024029198218e420000",
			INIT_37 => x"03e000088fb000108fb100148fb200188fb3001c8fb400208fb500248fb60028",
			INIT_38 => x"026028210c0000080200202100403021020020210c00001b8e50000427bd0030",
			INIT_39 => x"af82809c0800019c006210253042000f000519008f82809c00000000080001b5",
			INIT_3A => x"00808821afb100148c500000afb000100043102127bdffc82782801400041880",
			INIT_3B => x"afb40020afb50024afb60028afb7002cafbe0030afb3001cafbf003402002021",
			INIT_3C => x"122200bf24020001278580c10c0000080200202100403021afb200180c00001b",
			INIT_3D => x"8f8280a01622006a240200041222009e240200031222005124020002279380c0",
			INIT_3E => x"2795802c27968028347778402a0200043c03017d245e0bb0241000013c020000",
			INIT_3F => x"001080c0321000078c51000002d21021321200388f9080b02414001414400036"
		)
		port map(
			DIA => dmem_write_out, DIB => x"ffffffff",
			DOA => dmem_data_read, DOB => imem_data_out,
			ADDRA => dmem_addr(10 downto 2),	ADDRB => imem_addr(10 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_we, WEB => '0', DIPA => x"f", DIPB => x"f"
		);

	end generate; -- small_mem
	
	big_mem:
	if mem_type /= "small" generate
	begin
	
	dmem_data_ready <= '1';
	dmem_write_out <= dmem_data_in;
	dmem_bram_cs <= dmem_addr_strobe;
		
	dmem_0: RAMB16_S9_S9
		generic map(
			INIT_00 => x"0001210500000801fd00ff030006000801fb0001ff0000070000fa00c0019000",
			INIT_01 => x"f540f701422b8002421125203821c02121210800fa40214202012108210801fd",
			INIT_02 => x"802321c04023808010102f1d01245b1c03e0ac210800000242f125012300f302",
			INIT_03 => x"2f0a21107e2121241c202418d82008ac2121ffff1c04238023c0218021232300",
			INIT_04 => x"23002d2808181c202124f82bff0001000000218f240c2b00f503003001102121",
			INIT_05 => x"012150210b21141c18e0000801f7ff0100f70a305702010bff0108aa2101017a",
			INIT_06 => x"1801200814181cef2a230400e4b41c0d24042426b810b400042101fb40214202",
			INIT_07 => x"fc2a2304040c00fc2a2304040c080321023821004e102f14181ce09800200814",
			INIT_08 => x"00deb8b4d4a2049801fc2a23040013040c00fc2a23040013040c02080cef0100",
			INIT_09 => x"040c0821d4029404005102c0090414ff00000003022101c02101c3b4b00025a2",
			INIT_0A => x"082524b82000000300e0037b056100082121210080fc882304040c00fc882304",
			INIT_0B => x"de0007002008b4b01014181c00c00101e00100fc882304040c00fc882304040c",
			INIT_0C => x"218000009c25f09c2133211014181c20242c28d0213d80b4215d3f235d01c124",
			INIT_0D => x"081014181c2024282c08fa070d2421001521216823c0400183001412202121e8",
			INIT_0E => x"2024282c301c34212114001021c814809c9c250f009c00b521082121211b0430",
			INIT_0F => x"c007002138b014362c2840047db00100a06a049e035102c0bf01c1082121181b",
			INIT_10 => x"2121237326c32303000021082121284323211b2121002121082121144323211b",
			INIT_11 => x"8c8321b0803100c1040112142021218000011c0ab60044212e01212f21040308",
			INIT_12 => x"a08ca401210108002b0038081014181c2024282c3034b0f40ab60e8c4001b00e",
			INIT_13 => x"a08c02cdf4b6018c21a00421d640b6028ca034dedcb60c8ca034e5dcb6088ca4",
			INIT_14 => x"24282c303423c0ffb0a00e8c01a0a08c210ec3004db89b048ca000f134c8f4b6",
			INIT_15 => x"0000239bc0b0048c01048c21349823b6c0f4b0218c01218c2138b61014181c20",
			INIT_16 => x"b01814a8060501a80d242610b4b81412fc20141220e8141220d414121420c0e8",
			INIT_17 => x"726d69645066736320726d6961506f656b6d4120000000b4d0181421dda8b4d0",
			INIT_18 => x"206e7a6f206e636b6f447453725a6947006f4b655a6f696f5376560063656c20",
			INIT_19 => x"64087d589a501f48c9403734002c401cda1400ecdcc8b4000000006e676f7964",
			INIT_1A => x"000000000000000000000000000000000000000000008c0284047c0874026c04",
			INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(7 downto 0), DIB => x"ff",
			DOA => dmem_data_read(7 downto 0), DOB => imem_data_out(7 downto 0),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(0), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_1: RAMB16_S9_S9
		generic map(
			INIT_00 => x"0000180000000000ff00ff2e2e00000000ff0000ff0000000000ffe002008c00",
			INIT_01 => x"ff40ff0050104f003800280000182f4038100000ff20182800001800100000ff",
			INIT_02 => x"1828301931282918000000f300d9070000ff80100000000038ff28002000ff00",
			INIT_03 => x"000088000088800000000000ff0000801018ff7f000018181010181820201821",
			INIT_04 => x"20000000000000001000ff10ff0000000000180000001000ff2e2e0000002030",
			INIT_05 => x"0020c3880028000000ff000000ffff0021ff000000170000ff00000018000000",
			INIT_06 => x"00000000000000ff10100000008000001800101080808000008800ff28201800",
			INIT_07 => x"ff101000000000ff101000000000004000002820000000000000ff8000000000",
			INIT_08 => x"248080808000008000ff1010008800000000ff10100088000000000000ff0000",
			INIT_09 => x"000000100000000000000000000000f902040600008000804800108080002000",
			INIT_0A => x"003810800006001e1eff0000000000002830101910ff131000000000ff131000",
			INIT_0B => x"ff000006000080800000000000ff0000ff0000ff131000000000ff1310000000",
			INIT_0C => x"1010210080100080b000300000000000000000ff100100ff400100400100ff10",
			INIT_0D => x"00000000000000000000ff00001098000088908018101900100000000020a080",
			INIT_0E => x"00000000000000208800000010ff801880011000198000012800203020000000",
			INIT_0F => x"800000100080000080807800010b000080000000000000800000800020300000",
			INIT_10 => x"2028200020172081000028002030002828200080900010200030280028282000",
			INIT_11 => x"01282080200211ff000000000020202011000000000000100000280030000000",
			INIT_12 => x"8001800020000000020000000000000000000000000080ff0000000128008000",
			INIT_13 => x"800100ff0100000128800080ff1f0000018000ff050000018000ff0500000180",
			INIT_14 => x"0000000000202001808000010080800120002800000b0200018000ff00ff0100",
			INIT_15 => x"00002002208000010000012000ff200020018028010028012000000000000000",
			INIT_16 => x"80000080000000800010108080800000800000000080000000800000000080ff",
			INIT_17 => x"0061206a6f6f656e20006120726f726d6961756b000000800100002002808001",
			INIT_18 => x"206f65007a6f7200767500700061636f007661626164206e6c6175006920614e",
			INIT_19 => x"0c00020c010c010c000c000c000cff0cfe0c0c0b0b0b0b010000000072776500",
			INIT_1A => x"000000000000000000000000000000000000000000000c000c000c000c000c00",
			INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(15 downto 8), DIB => x"ff",
			DOA => dmem_data_read(15 downto 8), DOB => imem_data_out(15 downto 8),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(1), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_2: RAMB16_S9_S9
		generic map(
			INIT_00 => x"828400408200e084c085c60505c000e0a5c0a284c68200c00000001b001d9c1c",
			INIT_01 => x"a0084063058502e2076b2a0b00000500a060e0008004640540a2008060e06340",
			INIT_02 => x"05a2c30707a30202a7a600a5054402bf80bd8400e0c400c0076b2a08850040e2",
			INIT_03 => x"0005c0b20000a080b1b2bfb0bdbde08360624202bf6143034404620387866506",
			INIT_04 => x"04a202bde0b0b1b2c0bf40036362100502652000bf4011258005024226a24040",
			INIT_05 => x"620003008080b0bfb1bd00e0a568a663044042464704a568a763080000a5b000",
			INIT_06 => x"b102bde0b0b1bf40515062000084bf606440438284838264708062a005850340",
			INIT_07 => x"404443626368004044436263676609000706004402b040b1b2bfbd8200bde0b0",
			INIT_08 => x"0485828485006482024044436244026362004044436244026363036202a9a500",
			INIT_09 => x"63716200022c0231004022022b120f0e19180d0c11000b9f004a028788624400",
			INIT_0A => x"6344ee828d446203026240624062c34000e24309094042436263700040424362",
			INIT_0B => x"590058e2bde08788b0b1b2bf003229c6afa50040424362636b0040424362636c",
			INIT_0C => x"4406066282a24282a08080b0b1b2b3b4b5bfb6bd0000022002000202004202ee",
			INIT_0D => x"e0b0b1b2b3b4b5b6bf52353140c2914215006484620202420262060005804383",
			INIT_0E => x"b4b5b6b7beb3bf0080b150b043bd8204820062420582000060000040000050bd",
			INIT_0F => x"101051d21290144095967702035e10028222022202220293220285000040b200",
			INIT_10 => x"c040820044048385440365002040a505822000b0b251d020004065a505822000",
			INIT_11 => x"0005008510001040021000060564821010104004006202004042e00000640600",
			INIT_12 => x"82008343404205000062bde0b0b1b2b3b4b5b6b7bebf85400400a500050485a5",
			INIT_13 => x"840005400400100000841100400400050084bf400400050084bf400400050084",
			INIT_14 => x"b5b6b7bebf4404428482a5000485820000a502000004000500840011bf400400",
			INIT_15 => x"000004000484050004050000bf400400041084000004000000bd00b0b1b2b3b4",
			INIT_16 => x"80bdbf84408284844043a28382850600840506000584060005840600bf0584bd",
			INIT_17 => x"006673656c726d6952006673656b00612074746d0000008500bdbf0000808500",
			INIT_18 => x"72006c00750076006e62006c00640073006172006700427361726b00636b7461",
			INIT_19 => x"0000000000000000000000000000ff00ff000000000000000000000065006c00",
			INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(23 downto 16), DIB => x"ff",
			DOA => dmem_data_read(23 downto 16), DOB => imem_data_out(23 downto 16),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(2), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_3: RAMB16_S9_S9
		generic map(
			INIT_00 => x"80240010800003241ca0240000180003241ca024249000180000103c0c3c373c",
			INIT_01 => x"1000142400000030001001240800000000000300140000001030001000032414",
			INIT_02 => x"00000000000000008f270c343c343caf14278f0103ac0010001401350000102c",
			INIT_03 => x"0c24002708020004afafafaf272703af0000343c8f0400000000000000000000",
			INIT_04 => x"00a02427038f8f8f008f140224a026a2828002088f1002a214000024268f0002",
			INIT_05 => x"300034001000afafaf2700032414a0240010282424002410a024240800242408",
			INIT_06 => x"8f2427038f8f8f1400008f000caf8f1400100000af8f8f8f8f00301400000010",
			INIT_07 => x"1400008f8faf001400008f8fafaf2400242400343caf14afafaf278f0027038f",
			INIT_08 => x"0027978f270c8faf241400008f343c8faf001400008f343c8faf24af24142400",
			INIT_09 => x"8fafaf0024112411001429241124242424242424240024270030008f8f8f000c",
			INIT_0A => x"af0000af10308f00002410281428801100030000001428008f8faf001428008f",
			INIT_0B => x"140010302703afaf8f8f8f8f001525241424001428008f8faf001428008f8faf",
			INIT_0C => x"000000afaf00308f001000afafafafafafafaf270008241101082901082c2900",
			INIT_0D => x"038f8f8f8f8f8f8f8f2616261402028e2400002700000030008f240c24020027",
			INIT_0E => x"afafafafafafaf0200af8caf00272700af080030008f0008020c0200020c8e27",
			INIT_0F => x"00328c02328f24142727342a3c24243c8f162412241224271224270c0200af0c",
			INIT_10 => x"0300000c000000278e8e020c0200240002020c02028c02020c0002240002020c",
			INIT_11 => x"0c00008f000800102a260c2424020000002414240caf24001030020c008f240c",
			INIT_12 => x"af0caf2c002c240008af27038f8f8f8f8f8f8f8f8f8f8f10240c300c00248f30",
			INIT_13 => x"8f0c2414240c260c008f240014240c240c8f8f14240c240c8f8f14240c240c8f",
			INIT_14 => x"8f8f8f8f8f0000308f8f300c248faf0c003000000c2408240c8f00168f14240c",
			INIT_15 => x"00000208008f240c24240c008f14020c00248f000c24000c0027088f8f8f8f8f",
			INIT_16 => x"af278faf1028248f1000008f8f8f240c2724240c2427240c2427240caf242727",
			INIT_17 => x"006f656c7500612075006f656e76006673736f00000000af08278f0008afaf08",
			INIT_18 => x"6500650074006500697200690061007000636c007200726b76006f0065756e70",
			INIT_19 => x"0000000000000000000000000000ff00ff000000000000000000000065006c00",
			INIT_1A => x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1B => x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map(
			DIA => dmem_write_out(31 downto 24), DIB => x"ff",
			DOA => dmem_data_read(31 downto 24), DOB => imem_data_out(31 downto 24),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(3), WEB => '0', DIPA => "1", DIPB => "1"
		);
		
	end generate; -- big_mem
end Behavioral;
