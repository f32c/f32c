library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use work.boot_block_pack.all;

package boot_rom_mi32el is

constant boot_rom_mi32el : boot_block_type := (
x"10", x"80", x"1D", x"3C", x"03", x"00", x"00", x"08",
x"21", x"F8", x"00", x"00", x"E8", x"FF", x"BD", x"27",
x"03", x"00", x"02", x"24", x"14", x"00", x"BF", x"AF",
x"80", x"FB", x"02", x"AC", x"FE", x"FF", x"03", x"24",
x"F0", x"FF", x"03", x"AC", x"21", x"20", x"00", x"00",
x"56", x"00", x"00", x"0C", x"00", x"02", x"05", x"24",
x"0F", x"80", x"04", x"3C", x"0C", x"80", x"89", x"34",
x"F2", x"01", x"28", x"91", x"55", x"00", x"07", x"24",
x"00", x"00", x"2A", x"91", x"FF", x"FF", x"26", x"91",
x"03", x"00", x"25", x"91", x"21", x"00", x"07", x"15",
x"02", x"00", x"2B", x"91", x"F3", x"01", x"2C", x"91",
x"AA", x"00", x"0D", x"24", x"1D", x"00", x"8D", x"15",
x"00", x"72", x"0A", x"00", x"00", x"10", x"18", x"24",
x"21", x"78", x"C6", x"01", x"19", x"00", x"F8", x"15",
x"00", x"CA", x"05", x"00", x"21", x"F8", x"2B", x"03",
x"02", x"00", x"E2", x"2B", x"15", x"00", x"40", x"14",
x"00", x"1B", x"1F", x"00", x"00", x"02", x"04", x"24",
x"56", x"00", x"00", x"0C", x"00", x"FE", x"65", x"24",
x"10", x"00", x"04", x"3C", x"20", x"00", x"0C", x"3C",
x"01", x"00", x"89", x"24", x"20", x"00", x"0A", x"24",
x"43", x"33", x"0C", x"00", x"10", x"FF", x"06", x"A0",
x"2A", x"28", x"89", x"01", x"0F", x"00", x"A0", x"10",
x"00", x"00", x"00", x"00", x"01", x"FB", x"0B", x"80",
x"01", x"00", x"68", x"31", x"0B", x"00", x"00", x"11",
x"00", x"00", x"00", x"00", x"00", x"FB", x"07", x"80",
x"09", x"00", x"EA", x"14", x"FF", x"FF", x"8C", x"25",
x"01", x"00", x"8C", x"25", x"E3", x"00", x"00", x"0C",
x"00", x"00", x"00", x"00", x"76", x"00", x"00", x"0C",
x"00", x"00", x"00", x"00", x"40", x"00", x"00", x"08",
x"00", x"00", x"00", x"00", x"FF", x"FF", x"8C", x"25",
x"EC", x"FF", x"80", x"15", x"43", x"33", x"0C", x"00",
x"0F", x"80", x"0D", x"3C", x"00", x"80", x"A2", x"35",
x"21", x"08", x"40", x"00", x"00", x"80", x"04", x"3C",
x"10", x"00", x"05", x"3C", x"24", x"E8", x"44", x"00",
x"04", x"00", x"A0", x"13", x"00", x"40", x"02", x"24",
x"00", x"00", x"40", x"BC", x"FE", x"FF", x"40", x"14",
x"FC", x"FF", x"42", x"24", x"21", x"F8", x"00", x"00",
x"08", x"00", x"20", x"00", x"25", x"E8", x"A5", x"03",
x"14", x"00", x"BF", x"8F", x"08", x"00", x"E0", x"03",
x"18", x"00", x"BD", x"27", x"01", x"FB", x"02", x"80",
x"01", x"00", x"43", x"30", x"FD", x"FF", x"60", x"10",
x"00", x"00", x"00", x"00", x"00", x"FB", x"04", x"80",
x"08", x"00", x"E0", x"03", x"FF", x"00", x"82", x"30",
x"E0", x"FF", x"BD", x"27", x"14", x"00", x"B0", x"AF",
x"21", x"80", x"80", x"00", x"40", x"FB", x"04", x"24",
x"1C", x"00", x"BF", x"AF", x"18", x"00", x"B1", x"AF",
x"8D", x"01", x"00", x"0C", x"21", x"88", x"A0", x"00",
x"40", x"FB", x"04", x"24", x"86", x"01", x"00", x"0C",
x"0B", x"00", x"05", x"24", x"02", x"2C", x"10", x"00",
x"86", x"01", x"00", x"0C", x"40", x"FB", x"04", x"24",
x"02", x"2A", x"10", x"00", x"86", x"01", x"00", x"0C",
x"40", x"FB", x"04", x"24", x"21", x"28", x"00", x"02",
x"86", x"01", x"00", x"0C", x"40", x"FB", x"04", x"24",
x"40", x"FB", x"04", x"24", x"86", x"01", x"00", x"0C",
x"FF", x"00", x"05", x"24", x"1C", x"00", x"BF", x"8F",
x"14", x"00", x"B0", x"8F", x"0F", x"80", x"05", x"3C",
x"21", x"30", x"20", x"02", x"18", x"00", x"B1", x"8F",
x"40", x"FB", x"04", x"24", x"00", x"80", x"A5", x"34",
x"6A", x"01", x"00", x"08", x"20", x"00", x"BD", x"27",
x"C8", x"FF", x"BD", x"27", x"2C", x"00", x"B7", x"AF",
x"28", x"00", x"B6", x"AF", x"24", x"00", x"B5", x"AF",
x"20", x"00", x"B4", x"AF", x"1C", x"00", x"B3", x"AF",
x"34", x"00", x"BF", x"AF", x"30", x"00", x"BE", x"AF",
x"18", x"00", x"B2", x"AF", x"14", x"00", x"B1", x"AF",
x"10", x"00", x"B0", x"AF", x"91", x"00", x"13", x"24",
x"A1", x"00", x"14", x"24", x"B0", x"00", x"15", x"24",
x"B1", x"00", x"16", x"24", x"A0", x"00", x"17", x"24",
x"82", x"12", x"11", x"00", x"4F", x"00", x"00", x"0C",
x"10", x"FF", x"02", x"A0", x"39", x"00", x"53", x"10",
x"92", x"00", x"44", x"2C", x"0B", x"00", x"80", x"10",
x"81", x"00", x"05", x"24", x"28", x"00", x"45", x"10",
x"90", x"00", x"06", x"24", x"03", x"00", x"46", x"14",
x"80", x"00", x"07", x"24", x"86", x"00", x"00", x"08",
x"21", x"90", x"20", x"02", x"F3", x"FF", x"47", x"14",
x"82", x"12", x"11", x"00", x"AF", x"00", x"00", x"08",
x"04", x"00", x"1E", x"24", x"37", x"00", x"54", x"10",
x"A2", x"00", x"4D", x"2C", x"05", x"00", x"A0", x"11",
x"00", x"00", x"00", x"00", x"EA", x"FF", x"57", x"14",
x"21", x"F0", x"00", x"00", x"C5", x"00", x"00", x"08",
x"21", x"80", x"00", x"00", x"3F", x"00", x"55", x"10",
x"00", x"00", x"00", x"00", x"E4", x"FF", x"56", x"14",
x"34", x"00", x"BF", x"8F", x"21", x"10", x"20", x"02",
x"30", x"00", x"BE", x"8F", x"2C", x"00", x"B7", x"8F",
x"28", x"00", x"B6", x"8F", x"24", x"00", x"B5", x"8F",
x"20", x"00", x"B4", x"8F", x"1C", x"00", x"B3", x"8F",
x"18", x"00", x"B2", x"8F", x"14", x"00", x"B1", x"8F",
x"10", x"00", x"B0", x"8F", x"08", x"00", x"E0", x"03",
x"38", x"00", x"BD", x"27", x"4F", x"00", x"00", x"0C",
x"00", x"8A", x"11", x"00", x"FF", x"FF", x"DE", x"27",
x"FC", x"FF", x"C0", x"17", x"21", x"88", x"51", x"00",
x"87", x"00", x"00", x"08", x"82", x"12", x"11", x"00",
x"21", x"58", x"00", x"02", x"04", x"00", x"0C", x"24",
x"03", x"46", x"0B", x"00", x"01", x"FB", x"09", x"80",
x"04", x"00", x"2A", x"31", x"FD", x"FF", x"40", x"15",
x"00", x"00", x"00", x"00", x"00", x"FB", x"08", x"A0",
x"FF", x"FF", x"8C", x"25", x"F8", x"FF", x"80", x"15",
x"00", x"5A", x"0B", x"00", x"87", x"00", x"00", x"08",
x"82", x"12", x"11", x"00", x"86", x"00", x"00", x"08",
x"21", x"80", x"20", x"02", x"C0", x"FF", x"D2", x"13",
x"C2", x"77", x"10", x"00", x"21", x"80", x"10", x"02",
x"4F", x"00", x"00", x"0C", x"25", x"80", x"0E", x"02",
x"21", x"78", x"D1", x"03", x"00", x"00", x"E2", x"A1",
x"21", x"80", x"50", x"00", x"C5", x"00", x"00", x"08",
x"01", x"00", x"DE", x"27", x"21", x"80", x"00", x"00",
x"21", x"10", x"00", x"00", x"B4", x"FF", x"52", x"10",
x"21", x"18", x"51", x"00", x"C2", x"C7", x"10", x"00",
x"21", x"C8", x"10", x"02", x"00", x"00", x"65", x"80",
x"25", x"F8", x"38", x"03", x"01", x"FB", x"04", x"80",
x"04", x"00", x"86", x"30", x"FD", x"FF", x"C0", x"14",
x"00", x"00", x"00", x"00", x"00", x"FB", x"05", x"A0",
x"21", x"80", x"BF", x"00", x"D1", x"00", x"00", x"08",
x"01", x"00", x"42", x"24", x"95", x"01", x"00", x"0C",
x"21", x"20", x"20", x"02", x"87", x"00", x"00", x"08",
x"82", x"12", x"11", x"00", x"21", x"40", x"00", x"00",
x"21", x"30", x"00", x"00", x"21", x"10", x"00", x"00",
x"6D", x"33", x"0A", x"3C", x"3E", x"20", x"0B", x"3C",
x"00", x"08", x"0C", x"3C", x"01", x"00", x"0D", x"24",
x"03", x"00", x"0E", x"24", x"53", x"00", x"0F", x"24",
x"0D", x"00", x"18", x"24", x"21", x"C8", x"00", x"00",
x"0D", x"0A", x"43", x"25", x"01", x"FB", x"05", x"80",
x"04", x"00", x"A7", x"30", x"FD", x"FF", x"E0", x"14",
x"00", x"00", x"00", x"00", x"00", x"FB", x"03", x"A0",
x"03", x"1A", x"03", x"00", x"25", x"48", x"79", x"00",
x"04", x"00", x"20", x"15", x"00", x"00", x"00", x"00",
x"FF", x"FF", x"19", x"24", x"EF", x"00", x"00", x"08",
x"32", x"6C", x"63", x"25", x"F3", x"FF", x"60", x"14",
x"FF", x"00", x"05", x"24", x"FF", x"FF", x"03", x"24",
x"02", x"00", x"07", x"24", x"1B", x"00", x"61", x"04",
x"00", x"00", x"00", x"00", x"00", x"48", x"02", x"40",
x"24", x"C8", x"4C", x"00", x"02", x"00", x"20", x"13",
x"21", x"20", x"00", x"00", x"FF", x"00", x"04", x"24",
x"C3", x"CC", x"02", x"00", x"FF", x"00", x"49", x"30",
x"FF", x"00", x"39", x"33", x"2A", x"48", x"29", x"03",
x"03", x"00", x"20", x"11", x"00", x"00", x"00", x"00",
x"0F", x"01", x"00", x"08", x"0F", x"00", x"84", x"38",
x"F0", x"00", x"84", x"38", x"10", x"FF", x"04", x"A0",
x"01", x"FB", x"04", x"80", x"01", x"00", x"99", x"30",
x"EC", x"FF", x"20", x"13", x"00", x"00", x"00", x"00",
x"00", x"FB", x"04", x"80", x"13", x"00", x"61", x"04",
x"F6", x"FF", x"89", x"24", x"05", x"00", x"8F", x"14",
x"FF", x"FF", x"19", x"24", x"21", x"10", x"00", x"00",
x"21", x"18", x"00", x"00", x"0F", x"01", x"00", x"08",
x"03", x"22", x"06", x"00", x"4A", x"00", x"99", x"10",
x"00", x"00", x"00", x"00", x"CD", x"FF", x"98", x"10",
x"20", x"00", x"89", x"28", x"DD", x"FF", x"20", x"15",
x"21", x"10", x"00", x"00", x"01", x"FB", x"02", x"80",
x"04", x"00", x"42", x"30", x"FD", x"FF", x"40", x"14",
x"00", x"00", x"00", x"00", x"FF", x"00", x"00", x"08",
x"00", x"FB", x"04", x"A0", x"04", x"00", x"39", x"2D",
x"05", x"00", x"20", x"13", x"00", x"49", x"02", x"00",
x"FF", x"00", x"05", x"24", x"FF", x"FF", x"03", x"24",
x"01", x"01", x"00", x"08", x"02", x"00", x"07", x"24",
x"61", x"00", x"82", x"28", x"03", x"00", x"40", x"14",
x"D0", x"FF", x"82", x"24", x"38", x"01", x"00", x"08",
x"E0", x"FF", x"84", x"24", x"41", x"00", x"99", x"28",
x"03", x"00", x"20", x"17", x"25", x"10", x"49", x"00",
x"C9", x"FF", x"84", x"24", x"25", x"10", x"89", x"00",
x"01", x"00", x"63", x"24", x"15", x"00", x"6D", x"14",
x"F9", x"FF", x"59", x"24", x"03", x"00", x"24", x"2F",
x"0D", x"00", x"80", x"10", x"04", x"00", x"49", x"28",
x"00", x"F0", x"04", x"3C", x"00", x"10", x"05", x"3C",
x"24", x"E8", x"04", x"01", x"00", x"80", x"02", x"34",
x"00", x"00", x"40", x"BC", x"FE", x"FF", x"40", x"14",
x"FC", x"FF", x"42", x"24", x"21", x"F8", x"00", x"00",
x"08", x"00", x"00", x"01", x"21", x"E8", x"A5", x"03",
x"FF", x"00", x"00", x"08", x"21", x"10", x"00", x"00",
x"FD", x"FF", x"20", x"11", x"00", x"00", x"00", x"00",
x"21", x"28", x"42", x"00", x"4A", x"01", x"00", x"08",
x"05", x"00", x"A5", x"24", x"04", x"00", x"6E", x"14",
x"06", x"00", x"A9", x"28", x"21", x"10", x"42", x"00",
x"4A", x"01", x"00", x"08", x"21", x"38", x"E2", x"00",
x"A8", x"FF", x"20", x"15", x"00", x"00", x"00", x"00",
x"06", x"00", x"65", x"14", x"2A", x"C8", x"A3", x"00",
x"02", x"00", x"00", x"15", x"21", x"30", x"40", x"00",
x"21", x"40", x"40", x"00", x"FF", x"00", x"00", x"08",
x"21", x"28", x"60", x"00", x"9F", x"FF", x"20", x"13",
x"01", x"00", x"64", x"30", x"9D", x"FF", x"80", x"10",
x"2A", x"48", x"67", x"00", x"9B", x"FF", x"20", x"11",
x"00", x"00", x"00", x"00", x"00", x"00", x"C2", x"A0",
x"FF", x"00", x"00", x"08", x"01", x"00", x"C6", x"24",
x"08", x"00", x"E0", x"03", x"00", x"00", x"00", x"00",
x"19", x"00", x"C0", x"10", x"FF", x"00", x"02", x"24",
x"00", x"00", x"82", x"A0", x"00", x"00", x"8C", x"8C",
x"00", x"01", x"83", x"31", x"FD", x"FF", x"60", x"10",
x"21", x"50", x"00", x"00", x"FF", x"FF", x"C6", x"24",
x"FF", x"00", x"07", x"24", x"02", x"42", x"0A", x"00",
x"0D", x"00", x"C0", x"10", x"00", x"4E", x"0C", x"00",
x"00", x"00", x"87", x"A0", x"03", x"00", x"CB", x"30",
x"03", x"00", x"60", x"15", x"25", x"50", x"28", x"01",
x"00", x"00", x"AA", x"AC", x"04", x"00", x"A5", x"24",
x"00", x"00", x"8C", x"8C", x"00", x"01", x"8D", x"31",
x"FD", x"FF", x"A0", x"11", x"00", x"00", x"00", x"00",
x"73", x"01", x"00", x"08", x"FF", x"FF", x"C6", x"24",
x"25", x"20", x"28", x"01", x"00", x"00", x"A4", x"AC",
x"08", x"00", x"E0", x"03", x"00", x"00", x"00", x"00",
x"00", x"00", x"85", x"A0", x"00", x"00", x"82", x"8C",
x"00", x"01", x"43", x"30", x"FD", x"FF", x"60", x"10",
x"FF", x"00", x"42", x"30", x"08", x"00", x"E0", x"03",
x"00", x"00", x"00", x"00", x"80", x"00", x"02", x"24",
x"01", x"00", x"82", x"A0", x"00", x"00", x"83", x"8C",
x"00", x"01", x"65", x"30", x"FD", x"FF", x"A0", x"10",
x"00", x"00", x"00", x"00", x"08", x"00", x"E0", x"03",
x"00", x"00", x"00", x"00", x"E0", x"FF", x"BD", x"27",
x"14", x"00", x"B0", x"AF", x"1C", x"00", x"BF", x"AF",
x"18", x"00", x"B1", x"AF", x"21", x"80", x"80", x"00",
x"00", x"80", x"11", x"40", x"02", x"24", x"11", x"00",
x"E8", x"03", x"05", x"24", x"C0", x"01", x"00", x"0C",
x"FF", x"0F", x"84", x"30", x"42", x"2F", x"11", x"00",
x"21", x"20", x"40", x"00", x"EB", x"01", x"00", x"0C",
x"01", x"00", x"A5", x"24", x"21", x"88", x"40", x"00",
x"0F", x"00", x"02", x"3C", x"41", x"42", x"43", x"24",
x"2A", x"30", x"03", x"02", x"04", x"00", x"C0", x"14",
x"21", x"20", x"00", x"02", x"EB", x"01", x"00", x"0C",
x"0A", x"00", x"05", x"24", x"21", x"20", x"40", x"00",
x"80", x"22", x"04", x"00", x"EB", x"01", x"00", x"0C",
x"E8", x"03", x"05", x"24", x"80", x"22", x"02", x"00",
x"EB", x"01", x"00", x"0C", x"21", x"28", x"20", x"02",
x"0F", x"00", x"07", x"3C", x"41", x"42", x"E8", x"24",
x"2A", x"48", x"08", x"02", x"04", x"00", x"20", x"15",
x"01", x"00", x"4C", x"24", x"21", x"50", x"8C", x"01",
x"C0", x"58", x"0C", x"00", x"21", x"60", x"4B", x"01",
x"02", x"FB", x"0C", x"A4", x"1C", x"00", x"BF", x"8F",
x"18", x"00", x"B1", x"8F", x"14", x"00", x"B0", x"8F",
x"08", x"00", x"E0", x"03", x"20", x"00", x"BD", x"27",
x"21", x"10", x"00", x"00", x"07", x"00", x"A0", x"10",
x"01", x"00", x"A3", x"30", x"02", x"00", x"60", x"10",
x"00", x"00", x"00", x"00", x"21", x"10", x"44", x"00",
x"42", x"28", x"05", x"00", x"C1", x"01", x"00", x"08",
x"21", x"20", x"84", x"00", x"08", x"00", x"E0", x"03",
x"00", x"00", x"00", x"00", x"01", x"00", x"C2", x"30",
x"08", x"00", x"40", x"10", x"2B", x"50", x"05", x"00",
x"C3", x"1F", x"05", x"00", x"C3", x"3F", x"04", x"00",
x"26", x"28", x"A3", x"00", x"26", x"20", x"87", x"00",
x"23", x"28", x"A3", x"00", x"23", x"20", x"87", x"00",
x"2B", x"50", x"05", x"00", x"2B", x"40", x"A4", x"00",
x"0C", x"00", x"00", x"11", x"21", x"10", x"00", x"00",
x"0A", x"00", x"A0", x"18", x"00", x"00", x"00", x"00",
x"21", x"28", x"A5", x"00", x"D5", x"01", x"00", x"08",
x"21", x"50", x"4A", x"01", x"03", x"00", x"20", x"15",
x"00", x"00", x"00", x"00", x"23", x"20", x"85", x"00",
x"25", x"10", x"4A", x"00", x"42", x"50", x"0A", x"00",
x"42", x"28", x"05", x"00", x"F9", x"FF", x"40", x"15",
x"2B", x"48", x"85", x"00", x"02", x"00", x"C6", x"30",
x"02", x"00", x"C0", x"10", x"00", x"00", x"00", x"00",
x"21", x"10", x"80", x"00", x"08", x"00", x"E0", x"03",
x"00", x"00", x"00", x"00", x"CB", x"01", x"00", x"08",
x"21", x"30", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
x"00", x"00", x"00", x"00", x"00", x"00", x"00", x"00",
	others => (others => '0')
    );

end boot_rom_mi32el;
