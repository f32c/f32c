-- Copyright (c) 2015, Smart Energy Instruments Inc.
-- All rights reserved.  For details, see COPYING in the top level directory.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package config is
constant cfg_ddr_ck_cycle: natural := 1000; -- check is this value correct
end package;
