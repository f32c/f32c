--
-- Copyright 2008, 2010 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
--

-- $Id$

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Xilinx libraries
library UNISIM;
use UNISIM.VComponents.all;

entity bram is
	generic(
		mem_type: string := "big"
	);
	port(
		clk: in std_logic;
		imem_addr: in std_logic_vector(31 downto 2);
		imem_data_out: out std_logic_vector(31 downto 0);
		imem_addr_strobe: in std_logic;
		imem_data_ready: out std_logic;
		dmem_addr: in std_logic_vector(31 downto 2);
		dmem_data_in: in std_logic_vector(31 downto 0);
		dmem_data_out: out std_logic_vector(31 downto 0);
		dmem_byte_we: in std_logic_vector(3 downto 0);
		dmem_addr_strobe: in std_logic;
		dmem_data_ready: out std_logic
	);
end bram;

architecture Behavioral of bram is
	signal dmem_wait_cycle, dmem_must_wait, dmem_we: std_logic;
	signal dmem_data_read, dmem_write_out: std_logic_vector(31 downto 0);
	signal dmem_bram_cs: std_logic;
begin
	
	imem_data_ready <= '1';
	dmem_data_out <= dmem_data_read; -- shut up compiler errors
	
	-- 32-bit wide memory with wait state insertion on byte / half word writes
	small_mem:
	if mem_type = "small" generate
	begin
	
	dmem_data_ready <= not dmem_must_wait;
	
	-- We need a read followed by a write cycle if storing a byte or half a word, so
	-- insert a wait state in such cases
	dmem_must_wait <= '1' when dmem_wait_cycle = '0' and dmem_byte_we /= "0000" and
		dmem_byte_we /= "1111" and dmem_addr_strobe = '1' else '0';
	
	process(clk, dmem_must_wait)
	begin
		if rising_edge(clk) then
			if dmem_wait_cycle = '0' and dmem_must_wait = '1' then
				dmem_wait_cycle <= '1';
			else
				dmem_wait_cycle <= '0';
			end if;
		end if;
	end process;
	
	dmem_we <= '1' when dmem_byte_we /= "0000" and dmem_must_wait = '0' else '0';
	dmem_write_out(7 downto 0) <= dmem_data_in(7 downto 0) when
		dmem_byte_we(0) = '1' else dmem_data_read(7 downto 0);
	dmem_write_out(15 downto 8) <= dmem_data_in(15 downto 8) when
		dmem_byte_we(1) = '1' else dmem_data_read(15 downto 8);
	dmem_write_out(23 downto 16) <= dmem_data_in(23 downto 16) when
		dmem_byte_we(2) = '1' else dmem_data_read(23 downto 16);
	dmem_write_out(31 downto 24) <= dmem_data_in(31 downto 24) when
		dmem_byte_we(3) = '1' else dmem_data_read(31 downto 24);
	
	dmem_bram_cs <= dmem_addr_strobe;
	dmem: RAMB16_S36_S36
		generic map(
			INIT_00 => x"00000000000000001000fffa3c1be0000c0002b43c1d0001379c8c603c1c0000",
			INIT_01 => x"24a500011cc0fffba0a200002484000124c6ffff908200000000000018c00007",
			INIT_02 => x"1cc0fffda085000024c6ffff00052e0300052e0018c000060000000003e00008",
			INIT_03 => x"80820000248400010000182110400005808200000000000003e0000824840001",
			INIT_04 => x"1040000230a2000100001821108000080060102103e00008246300011440fffd",
			INIT_05 => x"00a038210060102103e00008000000001480fffa000420400064182100052842",
			INIT_06 => x"00073842106b0011012a2825240b0020080000380000182100052fc000004021",
			INIT_07 => x"10a0fff5000840401440fff724630001000550420085102b00024f8030e20002",
			INIT_08 => x"00073842146bfff1012a28253508000100852023000000001040fff32ce20002",
			INIT_09 => x"1480000327bdffe08f8480ac0100102103e00008acc400000000000010c00002",
			INIT_0A => x"8fa7001027a600100c00002f34a5f31d3c0500013444d9243c02075bafbf001c",
			INIT_0B => x"0005188000a2282300c33021000719c00007314000a328230002298000021880",
			INIT_0C => x"00441023000410c0006218210003188000872021008620230065182300062100",
			INIT_0D => x"00601021006218213442ffff3c027fff8fbf001c046100040043182300031880",
			INIT_0E => x"afb1001cafb20020afbf0024afb0001827bdffd827bd002003e00008af8380ac",
			INIT_0F => x"0c00002f2405000a00c0882127b200100800007e0200882100a0802104800024",
			INIT_10 => x"1480fff500052e0300022e0024420030262600018fa200100040202102403021",
			INIT_11 => x"8202000080650000022018210800008f8fbf00241040000c0211102ba2250000",
			INIT_12 => x"00c010218fbf00241440fff80203102b2463ffffa062000026100001a2050000",
			INIT_13 => x"00042023a0a200002402002d27bd002803e000088fb000188fb1001c8fb20020",
			INIT_14 => x"a0a7ffff2463000124080008080000aa0000182124a5000124b000010800007a",
			INIT_15 => x"000421001040fff72842000a24460030244700570004170224a500011068000b",
			INIT_16 => x"afb1001827bdffe00000000003e0000824a500011468fff7a0a6ffff24630001",
			INIT_17 => x"30620001000020213403c350000088211080000b00802821afb00014afbf001c",
			INIT_18 => x"8f700004008088213062000114a0fffb00052840008520210003184210400002",
			INIT_19 => x"00641824104000040043102400821026af8480b88f8380108f8280b48f640000",
			INIT_1A => x"0051102a005010238f620004000000000c0000e4af8480b48fbf001c1460000d",
			INIT_1B => x"8fb100182402000127bd002003e000088fb000148fb100188fbf001c1440ffef",
			INIT_1C => x"afb20008afb3000c27bdfff08f8280980000000027bd002003e000088fb00014",
			INIT_1D => x"240700022406003800002821344420003c02004eafb000001440002fafb10004",
			INIT_1E => x"0044102a004310238f6200048f630004af67000caf6600082409000300004021",
			INIT_1F => x"1440fffc0044102a004310238f6200048f630004af68000c000000001440fffc",
			INIT_20 => x"8f630004af63000c24030002af6200082402000c14a9ffef24a5000100000000",
			INIT_21 => x"af62000c000000001440fffc0044102a004310238f620004344488003c020013",
			INIT_22 => x"240200011440fffc0044102a004310238f620004344488003c0200138f630004",
			INIT_23 => x"279080c000004821304a0001000210c38f8780b48f8880b08f620000af828098",
			INIT_24 => x"240ef9ff2419020024180400240d0600240c00032412000200008821240b0001",
			INIT_25 => x"11320004000000001440005029220002240200c0112b000924130004240f0014",
			INIT_26 => x"8f6200048f630004af72000caf62000800001021240200d4112c000224020094",
			INIT_27 => x"004310238f6200048f630004af71000c000000001440fffc2842138800431023",
			INIT_28 => x"1140000800002821020230210043102100091900000910801440fffc28421388",
			INIT_29 => x"00031e0300021e002462ffe0104000032862007b144000052862006180c30000",
			INIT_2A => x"af6c000caf6300080082382500ee102430e20600108d0020304406008f620000",
			INIT_2B => x"8f630004af6b000c000000001440fffc28421388004310238f6200048f630004",
			INIT_2C => x"24c6000114afffe024a50001000000001440fffc28421388004310238f620004",
			INIT_2D => x"af8880b08fb000008fb100048fb200088fb3000c000000001533ffc025290001",
			INIT_2E => x"2902ffc100ee10241459ffdf000000001058000727bd001003e00008af8780b4",
			INIT_2F => x"240200801120ffb501024021080001542902003f01024023080001542c420001",
			INIT_30 => x"afb50024afbf002cafb6002827bdffd000000000000000000000102108000134",
			INIT_31 => x"00a0b0211080003300803021afb00010afb10014afb20018afb3001cafb40020",
			INIT_32 => x"004410210006108000062100af620000af82809c00a21025304200f08f82809c",
			INIT_33 => x"000210838f620000240600140c00001224050020028020210043a021278380e8",
			INIT_34 => x"2415001500008821006490212784806800621823000210c00002194030420001",
			INIT_35 => x"8fbf002c265200081635fffa263100071440000d02c21024029198218e420000",
			INIT_36 => x"03e000088fb000108fb100148fb200188fb3001c8fb400208fb500248fb60028",
			INIT_37 => x"026028210c0000080200202100403021020020210c00001b8e50000427bd0030",
			INIT_38 => x"af82809c08000194006210253042000f000519008f82809c00000000080001ad",
			INIT_39 => x"00808821afb100188c500000afb000140043102127bdffd02782801400041880",
			INIT_3A => x"00403021afb2001c0c00001bafb30020afb40024afb50028afbf002c02002021",
			INIT_3B => x"122200a724020002279580c01222009324020001278580c10c00000802002021",
			INIT_3C => x"0c00001224050020278480d48f8280a01622004d24020004122200b924020003",
			INIT_3D => x"0c0000122406001424050020240600140c00001224050020278480e824060014",
			INIT_3E => x"323100078c530000025410213234003824100014279280288f9180b0278480fc",
			INIT_3F => x"0040302102a5282124a500140005284302022823026020210c00001b001188c0"
		)
		port map(
			DIA => dmem_write_out, DIB => x"ffffffff",
			DOA => dmem_data_read, DOB => imem_data_out,
			ADDRA => dmem_addr(10 downto 2),	ADDRB => imem_addr(10 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_we, WEB => '0', DIPA => x"f", DIPB => x"f"
		);

	end generate; -- small_mem
	
	big_mem:
	if mem_type /= "small" generate
	begin
	
	dmem_data_ready <= '1';
	dmem_write_out <= dmem_data_in;
	dmem_bram_cs <= dmem_addr_strobe;
		
	dmem_0: RAMB16_S9_S9
		generic map(
			INIT_00 => x"0001210500000801fd00ff030006000801fb0001ff0000070000fa00b4016000",
			INIT_01 => x"f540f701422b8002421125203821c02121210800fa40214202012108210801fd",
			INIT_02 => x"802321c04023808010102f1d01245b1c03e0ac210800000242f125012300f302",
			INIT_03 => x"2f0a21107e2121241c202418d82008ac2121ffff1c04238023c0218021232300",
			INIT_04 => x"23002d2808181c202124f82bff0001000000218f240c2b00f503003001102121",
			INIT_05 => x"012150210b21141c18e0000801f7ff0100f70a305702010bff0108aa2101017a",
			INIT_06 => x"1801200814181cef2a230400e4b41c0d24042426b810b400042101fb40214202",
			INIT_07 => x"fc2a2304040c00fc2a2304040c080321023821004e002f04080cf09800200814",
			INIT_08 => x"c02101c3b4b0009801fc2a23040013040c00fc2a23040013040c02080cef0100",
			INIT_09 => x"2304040c00fc882304040c0821d4029404005002c0090414ff00000003022101",
			INIT_0A => x"040c00fc882304040c082524002000000300e0037b056100082121210080fc88",
			INIT_0B => x"80b521543f235401c124df00071008b4b00004080c00c00101e00100fc882304",
			INIT_0C => x"83001412202121e8218000009c25f09c2133211014181c20242c28d000002134",
			INIT_0D => x"21082121211b0430081014181c2024282c08fa070d2421001521216823c04001",
			INIT_0E => x"a702c09301c10821211c1b2024282c212118001421d014809c94250f009c00ad",
			INIT_0F => x"2121144323211bc0070021381428b0fc121420141220e8141220d4a04d04b903",
			INIT_10 => x"407d040308218000237326c32303000021212c21082121284323211b00210821",
			INIT_11 => x"2c000edcb60884a4a084a40121010830b614181c2024282c640044002401212f",
			INIT_12 => x"b6018421a00421e640b60284a02ceedcb60c84a064280021300814181c202428",
			INIT_13 => x"0484212cc423b6c0f4b0218401218421b8280484a000f12cd8f4b6a08402ddf4",
			INIT_14 => x"210ec3004d30b66414181c2024282c0e844001b00e848321b02328c0b0048401",
			INIT_15 => x"20e8141220d414121420c0e830b62314181c202428c0ff2cb0a00e8401a0a084",
			INIT_16 => x"000000b4c8181421d1a8b4c8b01814a8060501a80d242610b4b81412fc201412",
			INIT_17 => x"5a6f696f5376560063656c20726d69645066736320726d6961506f656b6d4120",
			INIT_18 => x"ac9884000000006e676f7964206e7a6f206e636b6f447453725a6947006f4b65",
			INIT_19 => x"00005c0254044c0844023c0434087d289a201f18c910370400fc40ecdae4d0bc"
		)
		port map(
			DIA => dmem_write_out(7 downto 0), DIB => x"ff",
			DOA => dmem_data_read(7 downto 0), DOB => imem_data_out(7 downto 0),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(0), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_1: RAMB16_S9_S9
		generic map(
			INIT_00 => x"0000180000000000ff00ff2e2e00000000ff0000ff0000000000ffe002008c00",
			INIT_01 => x"ff40ff0050104f003800280000182f4038100000ff20182800001800100000ff",
			INIT_02 => x"1828301931282918000000f300d9070000ff80100000000038ff28002000ff00",
			INIT_03 => x"000088000088800000000000ff0000801018ff7f000018181010181820201821",
			INIT_04 => x"20000000000000001000ff10ff0000000000180000001000ff2e2e0000002030",
			INIT_05 => x"0020c3880028000000ff000000ffff0021ff000000170000ff00000018000000",
			INIT_06 => x"00000000000000ff10100000008000001800101080808000008800ff28201800",
			INIT_07 => x"ff101000000000ff101000000000004000002820000000000000ff8000000000",
			INIT_08 => x"804800108080008000ff1010008800000000ff10100088000000000000ff0000",
			INIT_09 => x"1000000000ff131000000000100000000000000000000000f902040600008800",
			INIT_0A => x"000000ff1310000000003810060006001e1eff0000000000002830101910ff13",
			INIT_0B => x"00ff400100400100ff10ff0000000080800000000000ff0000ff0000ff131000",
			INIT_0C => x"100000000020a0801010210080100080b000300000000000000000ff00001001",
			INIT_0D => x"280020302000000000000000000000000000ff00001098000088908018101900",
			INIT_0E => x"000080000080002030000000000000208800000010ff80188001100019800001",
			INIT_0F => x"3028002828200088000010000080808000000000000080000000808000000000",
			INIT_10 => x"7801000000280b00200020172081000010888020002830008080200000900020",
			INIT_11 => x"0000000500000180800180002000000000000000000000000000000000003000",
			INIT_12 => x"00000128800080ff1f0000018000ff0500000180000200100000000000000000",
			INIT_13 => x"00012000ff20002001802801002801200b0200018000ff00ff0100800100ff01",
			INIT_14 => x"2000280000000000000000000000000001280080000128208020022080000100",
			INIT_15 => x"0080000000800000000080ff0000200000000000002001008080000100808001",
			INIT_16 => x"0000008001000020028080018000008000000080001010808080000080000000",
			INIT_17 => x"6164206e6c6175006920614e0061206a6f6f656e20006120726f726d6961756b",
			INIT_18 => x"0b0b0b010000000072776500206f65007a6f7200767500700061636f00766162",
			INIT_19 => x"00000c000c000c000c000c000c00020c010c010c000c000c000bff0bfe0b0b0b"
		)
		port map(
			DIA => dmem_write_out(15 downto 8), DIB => x"ff",
			DOA => dmem_data_read(15 downto 8), DOB => imem_data_out(15 downto 8),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(1), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_2: RAMB16_S9_S9
		generic map(
			INIT_00 => x"828400408200e084c085c60505c000e0a5c0a284c68200c00000001b001d9c1c",
			INIT_01 => x"a0084063058502e2076b2a0b00000500a060e0008004640540a2008060e06340",
			INIT_02 => x"05a2c30707a30202a7a600a5054402bf80bd8400e0c400c0076b2a08850040e2",
			INIT_03 => x"0005c0b20000a080b1b2bfb0bdbde08360624202bf6143034404620387866506",
			INIT_04 => x"04a202bde0b0b1b2c0bf40036362100502652000bf4011258005024226a24040",
			INIT_05 => x"620003008080b0bfb1bd00e0a568a663044042464704a568a763080000a5b000",
			INIT_06 => x"b102bde0b0b1bf40515062000084bf606440438284838264708062a005850340",
			INIT_07 => x"404443626368004044436263676609000706004402b040b1b2b3bd8200bde0b0",
			INIT_08 => x"90004a0287886282024044436244026362004044436244026363036202a9a500",
			INIT_09 => x"43626371004042436263726200022c0232004022022b130f0e19180d0c12000b",
			INIT_0A => x"636b0040424362636c6382eee28d446203026240624062c34000024309094042",
			INIT_0B => x"022002000202004202ee590058bde08788b0b1b2b3003329c6afa50040424362",
			INIT_0C => x"02620600058043834406066282a24282a08080b0b1b2b3b4b5bfb6bd00000000",
			INIT_0D => x"60000040000050bde0b0b1b2b3b4b5b6bf52353140c291421500648462020242",
			INIT_0E => x"220295220285000040b200b3b4b5bf0080b150b043bd82048200624205820000",
			INIT_0F => x"40a5a50502600011315354341092918400060506000584060005848222022202",
			INIT_10 => x"a50564060040840482004404838544235451826000b040101002600053510060",
			INIT_11 => x"bf0040040005008482008343404205bd00b0b1b2b3b4b5bf0462020040420000",
			INIT_12 => x"00100000841100400400050084bf40040005008404006200bde0b0b1b2b3b4b5",
			INIT_13 => x"050000bf40040004108400000400000004000500840011bf4004008400054004",
			INIT_14 => x"00a5020000bd0004b0b1b2b3b4b5bfa500050485a50005008504000484050004",
			INIT_15 => x"0584060005840600bf0584bdbd0044b0b1b2b3b4b50442bf8482a50004858200",
			INIT_16 => x"0000008500bdbf000080850080bdbf84408284844043a2838285060084050600",
			INIT_17 => x"6700427361726b00636b7461006673656c726d6952006673656b00612074746d",
			INIT_18 => x"000000000000000065006c0072006c00750076006e62006c0064007300617200",
			INIT_19 => x"0000000000000000000000000000000000000000000000000000ff00ff000000"
		)
		port map(
			DIA => dmem_write_out(23 downto 16), DIB => x"ff",
			DOA => dmem_data_read(23 downto 16), DOB => imem_data_out(23 downto 16),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(2), WEB => '0', DIPA => "1", DIPB => "1"
		);
	dmem_3: RAMB16_S9_S9
		generic map(
			INIT_00 => x"80240010800003241ca0240000180003241ca024249000180000103c0c3c373c",
			INIT_01 => x"1000142400000030001001240800000000000300140000001030001000032414",
			INIT_02 => x"00000000000000008f270c343c343caf14278f0103ac0010001401350000102c",
			INIT_03 => x"0c24002708020004afafafaf272703af0000343c8f0400000000000000000000",
			INIT_04 => x"00a02427038f8f8f008f140224a026a2828002088f1002a214000024268f0002",
			INIT_05 => x"300034001000afafaf2700032414a0240010282424002410a024240800242408",
			INIT_06 => x"8f2427038f8f8f1400008f000caf8f1400100000af8f8f8f8f00301400000010",
			INIT_07 => x"1400008f8faf001400008f8fafaf2400242400343caf14afafaf278f0027038f",
			INIT_08 => x"270030008f8f8faf241400008f343c8faf001400008f343c8faf24af24142400",
			INIT_09 => x"008f8faf001428008f8fafaf0024112411001429241124242424242424240024",
			INIT_0A => x"8faf001428008f8fafaf00003010308f00002410281428801100020000001428",
			INIT_0B => x"241101082901082c29001400102703afaf8f8f8f8f001525241424001428008f",
			INIT_0C => x"008f240c24020027000000afaf00308f001000afafafafafafafaf2700000008",
			INIT_0D => x"020c0200020c8e27038f8f8f8f8f8f8f8f2616261402028e2400002700000030",
			INIT_0E => x"1224271224270c0200af0cafafafaf0200af8caf00272700af080030008f0008",
			INIT_0F => x"0002240002020c00328c023224278f270c2424240c2427240c24278f16241224",
			INIT_10 => x"343c8f240c00243c000c000000278c8e000027020c0200260002020c8e020c02",
			INIT_11 => x"8f0010240c240c8faf0caf2c002c2427088f8f8f8f8f8f8f24af24001030000c",
			INIT_12 => x"0c260c008f240014240c240c8f8f14240c240c8f2408af0027038f8f8f8f8f8f",
			INIT_13 => x"240c008f14020c00248f000c24000c002408240c8f00168f14240c8f0c241424",
			INIT_14 => x"003000000c2708248f8f8f8f8f8f8f300c00248f300c00008f0208008f240c24",
			INIT_15 => x"2427240c2427240caf2427272708008f8f8f8f8f8f00308f8f8f300c248faf0c",
			INIT_16 => x"000000af08278f0008afaf08af278faf1028248f1000008f8f8f240c2724240c",
			INIT_17 => x"7200726b76006f0065756e70006f656c7500612075006f656e76006673736f00",
			INIT_18 => x"000000000000000065006c006500650074006500697200690061007000636c00",
			INIT_19 => x"0000000000000000000000000000000000000000000000000000ff00ff000000"
		)
		port map(
			DIA => dmem_write_out(31 downto 24), DIB => x"ff",
			DOA => dmem_data_read(31 downto 24), DOB => imem_data_out(31 downto 24),
			ADDRA => dmem_addr(12 downto 2),	ADDRB => imem_addr(12 downto 2),
			CLKA => not clk, CLKB => not clk, ENA => dmem_bram_cs, ENB => '1', SSRA => '0',
			SSRB => '0', WEA => dmem_byte_we(3), WEB => '0', DIPA => "1", DIPB => "1"
		);
		
	end generate; -- big_mem
end Behavioral;
