--
-- Copyright 2008, 2010, 2011 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--
--

-- $Id: bram.vhd 116 2011-03-28 12:43:12Z marko $

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library xp2;
use xp2.components.all;


entity bram is
	generic(
		C_mem_size: string
	);
	port(
		clk: in std_logic;
		imem_addr_strobe: in std_logic;
		imem_addr: in std_logic_vector(31 downto 2);
		imem_data_out: out std_logic_vector(31 downto 0);
		dmem_addr_strobe: in std_logic;
		dmem_write: in std_logic;
		dmem_byte_sel: in std_logic_vector(3 downto 0);
		dmem_addr: in std_logic_vector(31 downto 2);
		dmem_data_in: in std_logic_vector(31 downto 0);
		dmem_data_out: out std_logic_vector(31 downto 0)
	);
end bram;

architecture Behavioral of bram is
	signal dmem_data_read, dmem_write_out: std_logic_vector(31 downto 0);
	signal dmem_bram_cs: std_logic;
begin
	
	dmem_data_out <= dmem_data_read; -- shut up compiler errors
	dmem_write_out <= dmem_data_in;
	dmem_bram_cs <= dmem_addr_strobe;

	G_16k:
	if C_mem_size = "16k" generate
	ram_16_0: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x01A150220708A0D08A19004400025001E2A1FE3F0244001001080D40A8970A23A1A0010001400000",
		INITVAL_01 => "0x000000000000000000010A4D118200074590E2FB0225F0DE20070211E8590A610000310007010054",
		INITVAL_02 => "0x0000103A111A200000101A2000200B000411A000082100C0080161E1960A080E4118041180410030",
		INITVAL_03 => "0x0BAD10000012051022D0008080E00F0184C1608010203002C0002D602000020901A010000010DA10",
		INITVAL_04 => "0x180400180C1A21D020000020D020000020909A100000101C0101410064D1024D1002D103A111A20B",
		INITVAL_05 => "0x08A0C01203002401008401E1110C8406C810283400415110451821D0AAD100004002881004818048",
		INITVAL_06 => "0x0028010AAF00010000180104819E011984008C640180900601038480108009E890BE0F02280082A6",
		INITVAL_07 => "0x1406A03A90014100325003216020110220410040090CC110310024107A14080A8010050FE1000010",
		INITVAL_08 => "0x002411620112698008310E0AA00012100101A6F8070600BEEC0B013012000801E00C5F160210623D",
		INITVAL_09 => "0x1A260090CB0221C1E0110E008078A8038110201A0622A0084001A0414048012180521008A1002891",
		INITVAL_0a => "0x01008180BC0280C100401100411804118010820009EA1120101E2911A80F1028A062881221B02291",
		INITVAL_0b => "0x0E09F07C110224411808110C00804F0009F0A0900808D0861D088D201224008D209A201A81018841",
		INITVAL_0c => "0x1200C0AE7F02C0E122E702AEA1D0CC1D0EC090F100088090C008240080060620400090062F00E80F",
		INITVAL_0d => "0x1E2280BEF60001A09C1F01ED10380410082110881680E090080901C08040080810080C1A0EA0228E",
		INITVAL_0e => "0x03A14010080288C0301302A141B8B1182C41020801084032841A6511A44801E09058000100411818",
		INITVAL_0f => "0x1826A00004118041180011010096340AA50000761121E0C84F0BE500B400178D21E0500A4330E851",
		INITVAL_10 => "0x000F01B41C062A10AA051400B19A5D06C33022A118C1303A21006F11B4C1014CC016B0058AA1860C",
		INITVAL_11 => "0x050D80A0250A054000560E6B500E8203EF00A0561AC4F1DC1F024F80AA05100091564B0A0AB1A405",
		INITVAL_12 => "0x01E10100CD1B62F02421102400641D1A0400AA0500001046DC18044062210565108CDC07EC116212",
		INITVAL_13 => "0x0222119EFB02021184F319C320581B162411E8C00902801012108E10D6EE08080090C0090CC0C250",
		INITVAL_14 => "0x1806401084118040284F0AA05080050CE1F1E0F3020250804503E1F002021844F10A01082FF00801",
		INITVAL_15 => "0x08208010041181408260000CF096B40020F046120180309E2E000C216407002C009E4D00861070F1",
		INITVAL_16 => "0x090C00888801048182130804C1F8420B64004021040CF0200D19C2E0C025078ED050B4004360628C",
		INITVAL_17 => "0x000DB13E801AC0B1C2F1022211E0180301101C1105681182E001C0C08C1C1EA0010283182411E0C0",
		INITVAL_18 => "0x002181D0D017E8B08C0411600016FB1828109801026F0068051065001011032011E2010B466038FC",
		INITVAL_19 => "0x1088C0088C0086600CF605AA60D0850A005140B40AA8F016441FE4010A5F08894174881406116290",
		INITVAL_1a => "0x0A050000D019CF00AA000B40B08A611280F0166508E081904C1E0C0020C418080102CC0381C170F8",
		INITVAL_1b => "0x09800006011E8FE040861FEC0022B31187C03A060241802040090CC01841010180108C00840110C5",
		INITVAL_1c => "0x0204203E100226500C8710001024B31F0860602F0A2D30361E03C2600A0600C0F028060683602032",
		INITVAL_1d => "0x178280C2B01088C1881010240110040020808041010081180411804102C218482006810220803601",
		INITVAL_1e => "0x0A28F0D68106866106B400C820CA5100C17018FA0384009C3808608162F103EF11E02E002B807011",
		INITVAL_1f => "0x0005A016450B0F01607408A88020C410204198101008411804102C202E841188F102640A0620C0F8",
		INITVAL_20 => "0x0C2B001E8B00C080860402E001C254102C1180511988009041008101108008841188000805A11055",
		INITVAL_21 => "0x0E450112450AA00018DE1F0B11420B0C0011080E1A0810E015030800305002897002200680701201",
		INITVAL_22 => "0x0A6510A08302404056920465208011162BB03641076610603112218100481801401813080B100A06",
		INITVAL_23 => "0x0000000000000000001019CA2190AF1480812AA11325A0A0DE100440BC0E01C35152BF1AAE01C451"
	)
	port map (
		DIA0 => dmem_write_out(0), DIA1 => dmem_write_out(1),
		DIA2 => dmem_write_out(2), DIA3 => dmem_write_out(3),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(0), DOA1 => dmem_data_read(1),
		DOA2 => dmem_data_read(2), DOA3 => dmem_data_read(3),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(0), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(0), DOB1 => imem_data_out(1),
		DOB2 => imem_data_out(2), DOB3 => imem_data_out(3),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_1: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x01E00044C001C0F0002001C001E0001E0021FECF0402001E00000F00161000073000021182018000",
		INITVAL_01 => "0x000000000000000000000C6000600000400000F20000F01E60000621E02C0404E0BA06018001A000",
		INITVAL_02 => "0x142E2056201641A03C251641A0424301C0010610070201E2F501E2B0060000613066440885515680",
		INITVAL_03 => "0x054B2022E00802204410170050007E00402180510040816460144B0042A10404E16C21142E201621",
		INITVAL_04 => "0x08A50172011640B042A11C45B042A11C40401621142E201600038001C0B2000B2004B20562216400",
		INITVAL_05 => "0x0220500000024111C0010002002201002000201000200020101E02B000B2034111C4E50063306844",
		INITVAL_06 => "0x10400004FF02221118200401103E1F034000020000A0000012042111C20103E1F03000040111E002",
		INITVAL_07 => "0x06E1600A600602201E200002B05E22044550AC64088451229002410120200220E020821FE2102821",
		INITVAL_08 => "0x004401E4020043A0000005AC01A0210203018E27060401ACD60E07300A0E0C62E01C2F126F204660",
		INITVAL_09 => "0x044030603E00023160220A673006031862204200044600600000A3000250060270002300A2F00002",
		INITVAL_0a => "0x05A20022D1044320402E0C044088550AA620C4F307EF2000211E0020403F004F2040330042804002",
		INITVAL_0b => "0x0200F01E01044210222D04012040FF0220F002080160B0002B000B000000020B0016041602B02402",
		INITVAL_0c => "0x000110A6FF0400B044B3004FA160121E2B1024F201C20022120440B0161F0400016000004011E0BF",
		INITVAL_0d => "0x1E4821FEF001E200161F11E020421103C2C004100420103C20022210160B01620080B1000B30422B",
		INITVAL_0e => "0x0422103C20042110420000C220220200411024E100011040011200002C1E00000022010401102202",
		INITVAL_0f => "0x040001A01102222044D0020210242204420000770EE200845F05E2004A000AA50024200A42004460",
		INITVAL_10 => "0x0002301008004B2044021C00E1C0CE01C01004B20582F00262040A002A1200012000B0004F301800",
		INITVAL_11 => "0x002040403204024000440860200630180F20403300C2F038311A0F00440208004088300403301022",
		INITVAL_12 => "0x07E02026100044F04810024B100020030B1044020A0050AA020021000402004F001E030562404421",
		INITVAL_13 => "0x0444001EF305442008F4004020020404402082120420D0002102212004FF006010221204422184C0",
		INITVAL_14 => "0x022011C401022220043F04402040020442F1F0F1054C20602205E2F044A00003F04400044FF064A2",
		INITVAL_15 => "0x020E00401102221044040020C000200001F0022001A0105E0100E1204000020000400202072002F0",
		INITVAL_16 => "0x044230621C040110202B02220182B01E40000202020DF0421A01C01002000021000420000B000411",
		INITVAL_17 => "0x016601DE001E0820E412040221E0200402201E021C0101E0F00042502E2704020000000A40204012",
		INITVAL_18 => "0x004210023001E00002010221A000100E40000010000F800000000E010A2201C021E0E20020701EB6",
		INITVAL_19 => "0x00211044220660711090012100E0D204002020110201F0201303E030E02F0062000011080E2060F0",
		INITVAL_1a => "0x0402000011022110440004201022001402F020020441B084021FE4104044068B00042100202000F3",
		INITVAL_1b => "0x03A10000011E4F1080031FE40040220000600C2004E2804023066310440200421188030880002002",
		INITVAL_1c => "0x0402405E2000A021000003402040221E0100682F0C41200421040400A4800201C042000620002000",
		INITVAL_1d => "0x040050045210422020200241D02011000080200203C4002222044330643006A0A004020440005E00",
		INITVAL_1e => "0x1840F1C4020420C000200001001A201002001AFB044110322004410044B205EB21E811004C000020",
		INITVAL_1f => "0x0002100211002F1000110021B04222044F2044221A601022220442005A100240F0040D05004000C0",
		INITVAL_20 => "0x0043103E0000000002010420A048E0024820E2020C483064020042218402040020E0000420000022",
		INITVAL_21 => "0x02020022020440000211020001E0000002000002004001E00E000000400204203024410001001C12",
		INITVAL_22 => "0x120901200204000004F408424000B21E402044A00440004002004030042204623030200003200401",
		INITVAL_23 => "0x000000000000000000000E6320C40600C2604C020C460040670E4760CC240047700C6608C6208092"
	)
	port map (
		DIA0 => dmem_write_out(4), DIA1 => dmem_write_out(5),
		DIA2 => dmem_write_out(6), DIA3 => dmem_write_out(7),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(4), DOA1 => dmem_data_read(5),
		DOA2 => dmem_data_read(6), DOA3 => dmem_data_read(7),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(0), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(4), DOB1 => imem_data_out(5),
		DOB2 => imem_data_out(6), DOB3 => imem_data_out(7),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_2: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x01E001101001E0F0000001E001E00000008000C00000801E00000F00020000000010080028002000",
		INITVAL_01 => "0x000000000000000000001C6A00000000000000F80000001E00000000000F0000F01E00022001E000",
		INITVAL_02 => "0x000081020002000000000200000031000000C60000C001E02201E82062000003000000000001E600",
		INITVAL_03 => "0x000100000002400010100460200430000000C4200100805030000100000010010020000000000200",
		INITVAL_04 => "0x00000046000200100000010010000000001002000000801E4001E001E01000010010101020802000",
		INITVAL_05 => "0x0000101000000001E0000008000000000000000000000000001E0010001000000010F00000000000",
		INITVAL_06 => "0x00000000FF00000000000000001E0F00200000000020800000100001E00001E0F00200000001E008",
		INITVAL_07 => "0x00000000000000001E0001080102880000000000000001E01000000020000000F000001FE0000080",
		INITVAL_08 => "0x010201E008110230000005EF01E008000201E000000201E0F0000000040F0008101E0F000F000000",
		INITVAL_09 => "0x000000000F0000010080000200000010080100000102000000004000002001080010800048100088",
		INITVAL_0a => "0x01E0000010000700000F0000000000000000101001EF8100001E0880000F000F8000001100200088",
		INITVAL_0b => "0x0008F00037000000000F00000000FF0008F0000000201014810001A010A00001C002E00200100008",
		INITVAL_0c => "0x00400060FF00002010200000104E0000020000F80BE0000000000010020F0000002080010301E01F",
		INITVAL_0d => "0x1E0301E0F0044001040F060001000001E07000000000301E00000000020100200000100002000002",
		INITVAL_0e => "0x0000001E000000010000006000000800000010F00000000000060000060F00000000000000000000",
		INITVAL_0f => "0x000001E00000000000F000000010080000A19C00000800300F10002000CE0000000C8A1442000030",
		INITVAL_10 => "0x14400000000103011020038610204100200010380080F0003008000006000000008000000F000800",
		INITVAL_11 => "0x12000004000140019C0000000040001E0FE004000008F01E001E0F011020018E0000001040000060",
		INITVAL_12 => "0x01E00000000102101000000400000000040010A000860000000000001008000F001E000100011080",
		INITVAL_13 => "0x11020002F0106A0000F0000000000010008000000000F0000000000000FF00000000000000008040",
		INITVAL_14 => "0x000001E000000000005F1102000860000011F0F0106900B4001028F010320025F010A00101F00030",
		INITVAL_15 => "0x000F000000000000100900004000800000F000800080011E1000A0000000000000000000050000F0",
		INITVAL_16 => "0x000000000F000000000500000080501F000000080004F0000501E000000000000000000005000000",
		INITVAL_17 => "0x006000A0000A0000000000000000001008801E080A0001E0F00000000C0500000000000100000000",
		INITVAL_18 => "0x0100000060000000000000003000000A000000000000800000000000008000A00000F00000601EF0",
		INITVAL_19 => "0x00000000000000611EF601E000C058018A8014000000000000000000C00000000000000C0F00A0F0",
		INITVAL_1a => "0x1000219C0000000110CA00020000000C0000000000005000000060000000000F0000000000000000",
		INITVAL_1b => "0x0080700000010F01400003E720000800000000C010083000000000000000000001E0000000000008",
		INITVAL_1c => "0x000070028000E081E0000060000008020000E4000700800080000A00E0F000004000000E0000E000",
		INITVAL_1d => "0x100000000006000000800000F00000000030000001E0000000000000000000E0F000080000001E00",
		INITVAL_1e => "0x1F0011F00010007000800000000E001E080008F70000000E80010000108801E881F4000007000080",
		INITVAL_1f => "0x19400040000000000000000050000001030000001E000000000000000E00000010000711E0A00040",
		INITVAL_20 => "0x000500000000000000000000301000000800A0000003000008000001E000000800A0000100001008",
		INITVAL_21 => "0x0000A00008110A41C000000001E0000000000000000001E00F000001000010000000000000001E00",
		INITVAL_22 => "0x100801000000000000F800080000881F008000800000010000000000000000000010000005001020",
		INITVAL_23 => "0x000000000000000000101FEBA13C060E22F1426A180160807105E511C209012FC0061313C1012080"
	)
	port map (
		DIA0 => dmem_write_out(8), DIA1 => dmem_write_out(9),
		DIA2 => dmem_write_out(10), DIA3 => dmem_write_out(11),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(8), DOA1 => dmem_data_read(9),
		DOA2 => dmem_data_read(10), DOA3 => dmem_data_read(11),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(1), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(8), DOB1 => imem_data_out(9),
		DOB2 => imem_data_out(10), DOB3 => imem_data_out(11),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_3: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x01E080240011E0F0103001E801E08800002000C00602401E00100F010000000000000F0004000080",
		INITVAL_01 => "0x0000000000000000000006C000000000800000FC0000001E00000040001F0200F01E00080001E008",
		INITVAL_02 => "0x0100404020004801003000480050200000000400100201E00801E20040000000000000000001F400",
		INITVAL_03 => "0x1800211000000FA1220000408000200000000080010890042001000050080E000000280100600028",
		INITVAL_04 => "0x00000004000040005008008000500800600000280100101E0001E001E00200002004020402200400",
		INITVAL_05 => "0x1100001E00110001E0080004011008010000000800008000001E0200000210080002F00000000000",
		INITVAL_06 => "0x00200002FF11018000100000001E8F00080010000000F00088100001E00001E8F10000080881E002",
		INITVAL_07 => "0x0000000000000B001E0001E20160981120000000000001E00000400000800000F100011FE1810028",
		INITVAL_08 => "0x016001E6021F6020000001EF01E0B5000001E000000001E0F0000000000F0002001E0F000FB00000",
		INITVAL_09 => "0x002000000F0006000022000000000000022120000D40000000000000000001E2001E2000090000F2",
		INITVAL_0a => "0x01E0000000060000000F0000000000000010160001EF21E0C01E0F20000F004F70E0001E4B0020F2",
		INITVAL_0b => "0x000FF00002130000000F00000000FF000FF0100000000004200000201E2010002000200008000008",
		INITVAL_0c => "0x00000000FF1004000400000000100000000010F213E0000000002000008F02000000F0010081E00F",
		INITVAL_0d => "0x1E2081E0F0000200400F000091000001E81010000200001E00000100000000080000000080010080",
		INITVAL_0e => "0x0608001E000200002000000300000801000002F00000002000000000000F00000000000000000008",
		INITVAL_0f => "0x100001E00000000000F000010018C70EC5608600000C00820F1807C0C05400000006211400000000",
		INITVAL_10 => "0x020000000000402134C9010700000000000012020001F0000200000000020000800000010F000000",
		INITVAL_11 => "0x140001420419EA00EC0000004040001E0F306200000FF01E001E0F0110A700C500000010A0000034",
		INITVAL_12 => "0x11E000100001060098C00080000090008000B42B01410000000000001206004F000000040000943B",
		INITVAL_13 => "0x04A60000F004049012F0000000000005008000000000F0001400001006FF00000000000000000200",
		INITVAL_14 => "0x000001E000000000020F0D26200A4000080004F00401100400020FF0040C0020001EC000E0F00002",
		INITVAL_15 => "0x000F000000000100180700000000600000F000200000009E40000000E000000000000000008000F0",
		INITVAL_16 => "0x000000000F000000001000000000001EA00000020000F0400001E000000000000000200000001000",
		INITVAL_17 => "0x0040000000000060000000000000400203201E01000001E0F0000000002000000000000100800000",
		INITVAL_18 => "0x00840000000000000000000000000000400000000000700000000000208000002000F20000001EF0",
		INITVAL_19 => "0x00000000000000003EF001E000000B0E86500600000000000000000000000000000000000F2000F0",
		INITVAL_1a => "0x0803504200000001F8670C05000000000000000000000000000000010000000F0002800000800000",
		INITVAL_1b => "0x000000000000CF00A00001E00120430000000010100A012000000000000A000801E0000000000005",
		INITVAL_1c => "0x0A00006050000011E0000000F1E01F0000001E000040900E6006090006F000000040000000000000",
		INITVAL_1d => "0x020000120000000000800100F00000000000000801E000000000000002000000F0120F1940009E00",
		INITVAL_1e => "0x1EA001E803100000001000000000401E020000F00E00000080086000740205E021F20000E0000080",
		INITVAL_1f => "0x0AC50080000000000000000000400000400000801E0000000000200020000000000E0005E0600000",
		INITVAL_20 => "0x00400000000000000000080000000001202000090000000008000801E000000020000000000000C7",
		INITVAL_21 => "0x000290000F0ECC608000000001E0000000000000000001E00F000000E00018000012000000001E04",
		INITVAL_22 => "0x000000000102000008F20A245000021E8030AA0002A0004002002000000000010000900000200630",
		INITVAL_23 => "0x000000000000000000000E63204C070847606C600C4660C063064660CC7600C5600C650CC670C003"
	)
	port map (
		DIA0 => dmem_write_out(12), DIA1 => dmem_write_out(13),
		DIA2 => dmem_write_out(14), DIA3 => dmem_write_out(15),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(12), DOA1 => dmem_data_read(13),
		DOA2 => dmem_data_read(14), DOA3 => dmem_data_read(15),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(1), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(12), DOB1 => imem_data_out(13),
		DOB2 => imem_data_out(14), DOB3 => imem_data_out(15),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_4: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x000840000013A000A40C00E90010640880807026000B2000580A004130081FCDC0F6A000000064D0",
		INITVAL_01 => "0x0000000000000000000001E6300C2000A04012550B20810C001EA0409C8410094004020400002074",
		INITVAL_02 => "0x174A000005000880EE0500022006401A60600A450A00E00A041C000080E400001046450CEEF1B80C",
		INITVAL_03 => "0x04A000A42000E0000000008F3088400AE0700C540C030000420A005002100000000A0E1DAD00A00B",
		INITVAL_04 => "0x0FCF0008C500050016BA14050010870E0000A002048400529008C100E6000A4000A0000000000050",
		INITVAL_05 => "0x0860000000040F01A00B0D67A100070B80C0A846000321A0F500A000AA000882F040DD0001206856",
		INITVAL_06 => "0x0C030004030CA270CE031A0011E4201E01000403000000002001E011BA001E4701402A0727200C03",
		INITVAL_07 => "0x0EA0604A5315204044240E00000000000450DCF0024371BA05000F5008021E02D0A052006280EE56",
		INITVAL_08 => "0x0800600E4000C060680200C0D1863012C040AA221E6041DC991E0851804F1FC0008847008A0010E0",
		INITVAL_09 => "0x08CDD060301C609016001760A0124C0060001C53180031008C1807706606080040E0040E0000E800",
		INITVAL_0a => "0x03AD01EE0F00E570CA5D1A001046450CEE01F203126000083406E0008A530000E0EE22000500CE00",
		INITVAL_0b => "0x0000100601000F00243D1A0011E00104401008030801008200088000000004800080050080001E40",
		INITVAL_0c => "0x06A4F00801000500800402005008F00020F0042009AD0002231E0400803000024000000040406802",
		INITVAL_0d => "0x06005000000A000040430001001E0105A22004D005E001FAD00020F08040080000880F00A0400030",
		INITVAL_0e => "0x0080F01AD00001F002300E00509E000A0F0020D2000DF0040F00402080FD00A62006001A00105E23",
		INITVAL_0f => "0x00E0610601046450DED21A0001F0641B69010A0B10A060C82411EDF17AA81F4890EA240E44900A07",
		INITVAL_10 => "0x1EE2F04029120001086109E361E40301A9C180001E0000A8000040B00000000400040A1409904000",
		INITVAL_11 => "0x04A200C66F0D2F61D89E1860B156A20122610683040590A0550106109E2D1F85218A500924904E82",
		INITVAL_12 => "0x066D0016B2018441F00F1D8021FE320180A0AE940EC390C62007CDC1C8C3164AB00A200A0F00AC40",
		INITVAL_13 => "0x1A8221A8201402114222050870EC2006030000231E22D000400E8700042507A00024340ACFF00003",
		INITVAL_14 => "0x1E0111BA000243F05E0F1962A1727212E661C2200401600462022120120113E020068111CE200600",
		INITVAL_15 => "0x004D51A00105E0F1FE1210450040CC084BB0400A0008010E16100F00AA4008858004200640000412",
		INITVAL_16 => "0x08A671E01D1A0011E4001A4D501E02014A9040800280100020000C700AC60CA7004033024000401F",
		INITVAL_17 => "0x1B00800650004080B63B04E090D67A0100009E3001E71062270CA430000004065002040803006423",
		INITVAL_18 => "0x17ADF0FC0001A76040541E05008E020002F1F22A1503311CDD1D8C91607B0A0650C62501E2010CE0",
		INITVAL_19 => "0x00012068560FE2007490060F200E0E096C808CC80C40505E9F014870040203E00060FF0080001ACC",
		INITVAL_1a => "0x11A570827C1081F130CE1709E17288004060A8200E0400A603020450005F002D000050000020404D",
		INITVAL_1b => "0x0A020000F01D8CE1283014E06000260CA100802200000000360FCF104A50088001BA0003EDC000BA",
		INITVAL_1c => "0x172700880502032042300A0400002912661006070004E01AEC1C02600A54100F000AF1004740000E",
		INITVAL_1d => "0x02822040030085F04A040200D1A00F000001E85001AD00022308A671C0F11E0901FC8E1DC9F17C9B",
		INITVAL_1e => "0x002AC0026306A200A0440440F100720E60408040000550A088086500400000800086030A00000800",
		INITVAL_1f => "0x1589E0F8970406509203000200045F0000F08A001BA00024340A0F2000E913E081FA50022210080B",
		INITVAL_20 => "0x0000A00E65008031004300040080380400000400006041E450082001BA001E00001EF91E020100FE",
		INITVAL_21 => "0x0A842084F91D88A11C8A10E760865708A430C833044F31D0981BEC813CDC0163014000132A000050",
		INITVAL_22 => "0x00C0600009000000CA0514AAA000050000214A0404A340A0100003D000120680F00001020000F65B",
		INITVAL_23 => "0x00000000000000000000016CB00A0F1F452008F00AC4F0001E06AB40282A01AE8002240624214C00"
	)
	port map (
		DIA0 => dmem_write_out(16), DIA1 => dmem_write_out(17),
		DIA2 => dmem_write_out(18), DIA3 => dmem_write_out(19),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(16), DOA1 => dmem_data_read(17),
		DOA2 => dmem_data_read(18), DOA3 => dmem_data_read(19),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(2), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(16), DOB1 => imem_data_out(17),
		DOB2 => imem_data_out(18), DOB3 => imem_data_out(19),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_5: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x00080000200240A080020041001800198A6048000104001400000820280100000000000044608010",
		INITVAL_01 => "0x0000000000000000000004466018C000C8604E2000E040E8000C00808C8808498010480040014080",
		INITVAL_02 => "0x0040000000000C01800000080008A000040014A0100000800800800180000960B176BB176BB17201",
		INITVAL_03 => "0x1A00013000002300000001C191E2A00164A0008A02011000410200001E1F00001000080100000002",
		INITVAL_04 => "0x176B0010000000000402000000180C000000000600C0002211146300AE000CA000C0000000000060",
		INITVAL_05 => "0x1100000804110BB160E80480E110E8190E00180000C4017CB014800000000C06B000BB1D6BB176BB",
		INITVAL_06 => "0x140001D466110480000017CBB160801601009064000040088A116BB176EB1608C100021CC8819408",
		INITVAL_07 => "0x0C2C60AC04000010B0041E028000EC150BB176BB176BB17600160B0000881760B11C000CC48118A8",
		INITVAL_08 => "0x0D80D11AC201E0702EC501AA80C86018E040C0600E0040E271020770C04600C2008C010C26000C0E",
		INITVAL_09 => "0x01E80174A41AE4A018240880A1144A014680161000000150660C0A600001020201E0200C0801EE02",
		INITVAL_0a => "0x176BE1740B014AA140AB17CBB176BB176BE17E0B16E620009B0FE0201217150EC0BEAA004701FE02",
		INITVAL_0b => "0x0408310201150BB176BB17CBB160231548311064000100020000001008141000100012000A017608",
		INITVAL_0c => "0x0000B00023088000000002050000B00B60B17000016BE176BB160000008406200000600C2080A000",
		INITVAL_0d => "0x0000800214000241600001E4C156BB176801D0BE01600176BE1760B00000000880800B0800008880",
		INITVAL_0e => "0x1508B176BE0D6BB0020400020116AA090BB160B801CBB000EB00044100BB018800D00817CBB17608",
		INITVAL_0f => "0x128C00C8BB176BB176B817C2B162EC108E100010000060840E1A2800400000001180600000108000",
		INITVAL_10 => "0x020010080502C0016A1D020110000114014000001600A0800000064000000100900008092E0000B0",
		INITVAL_11 => "0x0260808001122A100010000080000105CF00800001C2B0140101AB10781600001000120800001806",
		INITVAL_12 => "0x13660010000440006209110010C0D00800015805000000000402C0000E4B1080014804020B203EB0",
		INITVAL_13 => "0x1001500804040151020C1180C0100A1508A096BB176AB01C00150801946A116EB176BB176BB00001",
		INITVAL_14 => "0x1769B176EB176BB0140C0D010000010000A002040C01A0006603E30082011220E046131E04008E00",
		INITVAL_15 => "0x160B817CBB176010601102000014A8000A000844000121D818020BC0500A00C01086061000805652",
		INITVAL_16 => "0x176BB176BB17CBB1600000020016000C820000440A00105C20010221442A0042A010A212008150BB",
		INITVAL_17 => "0x0186100C000008B1B8DC1BC2C0C020002000EC6E01C131E6F20221100000038A20060401448014BB",
		INITVAL_18 => "0x018801600015CC801480008000024E0004302E4000EE00E0E00040E0142C1408E08CCE1C600014CA",
		INITVAL_19 => "0x1D6BB176BB17600000D00DCC0002021400E04022040A41C61B0807B000430F6511C8000004001462",
		INITVAL_1a => "0x19060002EA1DCF117E0009E0E1DC02000CA11C0E148A01544A1A0AA110AB176B01C08A148480108B",
		INITVAL_1b => "0x000000040C16CC900014042011C0FA0001808C00088E019CBB176BB1760A1168B176EB1760000002",
		INITVAL_1c => "0x100C014C0002002002040000E088FD0E2010024601009190700AC1001000168A01C00100050000C4",
		INITVAL_1d => "0x120140084B016BB160A8170BB17CBB0080017008176BE176BB176BB164B11600416A131F2B01CE46",
		INITVAL_1e => "0x10A0204E0B0601002CA4002E500061002450001001400000201E20C14806112060428B0000004286",
		INITVAL_1f => "0x0000600C66018A80C26002800014AB0800B1548B176EB176BB168B10800D0360F008000A21108000",
		INITVAL_20 => "0x080001D8A60120901060088000201000800014240960B1760A1168B176EB1620000231160050206A",
		INITVAL_21 => "0x0C4700EC3F1441000C760C46C0EC66158060CE711C07604E3100E0F0E00000024000000000001404",
		INITVAL_22 => "0x00000000E00500C18840008200000A140EA0800800040000A00D0CB1D6BB1764B0004502C0005806",
		INITVAL_23 => "0x0000000000000000000000A3200E060C06704C500CC65040220EE670CC7600C7700C740CC670C000"
	)
	port map (
		DIA0 => dmem_write_out(20), DIA1 => dmem_write_out(21),
		DIA2 => dmem_write_out(22), DIA3 => dmem_write_out(23),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(20), DOA1 => dmem_data_read(21),
		DOA2 => dmem_data_read(22), DOA3 => dmem_data_read(23),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(2), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(20), DOB1 => imem_data_out(21),
		DOB2 => imem_data_out(22), DOB3 => imem_data_out(23),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_6: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x00200000D800E04000030060002000110400600400000008150004300A8408844098C011A00198C0",
		INITVAL_01 => "0x0000000000000000000001834108000204806070120100808008A800080400E841084801A8008040",
		INITVAL_02 => "0x082400180418004008041800400058188041887C0F80C088C71880C0B0C401ECF1FEFF1FEFF0EE8C",
		INITVAL_03 => "0x068C004440188200008018EC70484819E0718877080001846C080C400241000C4188010824009801",
		INITVAL_04 => "0x1FEF018AC41804C002410804C000400800C098000804018C460EC600CCC004CC0040C00180018027",
		INITVAL_05 => "0x0660C000001E0FF0E033022140E6330863408840000000E6F40800C088C00080F0807707EFF1FEFF",
		INITVAL_06 => "0x000400604401800088040E6FF1E8F61F0000864001800000F001EFF0EE3F1E870070110087F09820",
		INITVAL_07 => "0x1880C0C042088040C8420C42001000000FF1FEFF1FEFF0EE841E4F4188041FE47006410880C00800",
		INITVAL_08 => "0x1C086084220448618C6610C1D0841005C82088040088208804086C01D02408028048440080003840",
		INITVAL_09 => "0x084641E4F40EC0F186110888F01E8F19E0100E44000841EA6E1D0F608884084240C4240D0280CC22",
		INITVAL_0a => "0x1EE731FECF00E4F1F8F70E6FF1FEFF1FEF21E48F1EC62046270CC22084460445200CFF0442804C22",
		INITVAL_0b => "0x0400600884000FF1FEF70E6FF1E0661FE0601E000984C0802C088C0000001E8C0098061880C1FE40",
		INITVAL_0c => "0x0884F10866000CC080C418C04188F601ECF1FE4008E731FEFF1E04C098FC04C24180000048F088C4",
		INITVAL_0d => "0x0808F0C46409824018441004001EFF1EEF007E7301E0C1EE731FE2F0984C098F4008CF098C4008FC",
		INITVAL_0e => "0x0000F1EE7301EFF01C440982601E00000FF1E07C0067F0083F10800018F700844000000E6FF1FE4F",
		INITVAL_0f => "0x1E04D080FF1FEFF1FE7C0E63F1E011022000002204400086C7038100240004424098000842408CC4",
		INITVAL_10 => "0x0082208840084C20440104002048820A444080C01F004004C210850058200082F1085C09E44090C6",
		INITVAL_11 => "0x0044200023040120002204450004260A00C0002208E340402207C6E04201040020442602022088C0",
		INITVAL_12 => "0x0E2521CE240C405060010228E0A8240408E0440004002044461CAEE084420824409840038F502020",
		INITVAL_13 => "0x024061C44403802180441804008040000C009EFF1FEC700610018000004418E3F1FEFF1FEFF10086",
		INITVAL_14 => "0x1FE4F0EE3F1FEFF0828504001040020442018044018001000004624086C0180830460202424082C2",
		INITVAL_15 => "0x1E87C0E6FF1FE0E0E6601DCEC0820C1C80408A0C018E5008001D0F1048E41C8EE0C440188800DE06",
		INITVAL_16 => "0x1FEFF1FEF70E6FF1E8081DC6E19E840A0DE08AC001CC4048E81C26209C64084240800E18884080FF",
		INITVAL_17 => "0x02C5410040108100180C0085C02224008000084210CE600C02188441D02C080C21CCE408000080FF",
		INITVAL_18 => "0x0220E03C800A0000800E1C8EC1C84218443080430801000E2408A420002C090020084207E480AA41",
		INITVAL_19 => "0x07EFF1FEFF1FE480064808AD411C81020000603306800066EF0A60F1082201E44020EE11C0218A11",
		INITVAL_1a => "0x00A000000F0000E02200020000002210840000401E87C1FE4701877018FF1FE70060F00804F08807",
		INITVAL_1b => "0x1D8E800AE70227001CE50288400A001DC40008C20080C018FF1FEFF1FE6019E0F0EE3F1FE6E1DCE1",
		INITVAL_1c => "0x042480000E09022084E01D8E30403205CE210002184310A22300402100421E8FC03CE211C421001C",
		INITVAL_1d => "0x01C440404F19EFF1EC0C1E0F70E6FF1C00C1F8601EE731FEFF1FEFF1E4F41F0E61C4E3024EE00A15",
		INITVAL_1e => "0x022E20A4E205C281C80C1C47C05024084041D848000EE1D02E000E4040C204CC20C0201C08E0DC04",
		INITVAL_1f => "0x00010000000800001C0E088EC04EFF084CF0FE0F0EE3F1FEFF1E4F4050E51DE311C0280482009CCE",
		INITVAL_20 => "0x084CE00000000000800E008EC090441C08218E6009ECF1FE6019E0F0EE3F1E88218C7E1F0401D011",
		INITVAL_21 => "0x02C20022E102200002110241408801000440A804068140E074062310284401C611C25E028E1008E0",
		INITVAL_22 => "0x10884100300200400050000100A080180000208800044000400000707EFF1FE2F1D004080C20C001",
		INITVAL_23 => "0x0000000000000000000001ADC01801080140702008282000A91F81F014F500E1200240040AF0A880"
	)
	port map (
		DIA0 => dmem_write_out(24), DIA1 => dmem_write_out(25),
		DIA2 => dmem_write_out(26), DIA3 => dmem_write_out(27),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(24), DOA1 => dmem_data_read(25),
		DOA2 => dmem_data_read(26), DOA3 => dmem_data_read(27),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(3), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(24), DOB1 => imem_data_out(25),
		DOB2 => imem_data_out(26), DOB3 => imem_data_out(27),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	ram_16_7: DP16KB
	generic map (
		-- CSDECODE_B => "000", CSDECODE_A => "000",
		WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
		GSR => "ENABLED", RESETMODE => "SYNC", 
		REGMODE_B => "NOREG", REGMODE_A => "NOREG",
		DATA_WIDTH_B => 4, DATA_WIDTH_A => 4,
		INITVAL_00 => "0x00238000A01420107001002800268A06610066020020400282140131040204422046300140110630",
		INITVAL_01 => "0x0000000000000000000000C32004A002012026200661302600024000620200222004120140000018",
		INITVAL_02 => "0x0542000002000A214402000A2014200641200423040030240206200040320B40A154AA154AA04603",
		INITVAL_03 => "0x0040015420004000000000432024200701200422040A000023040020142A000020040A054200400A",
		INITVAL_04 => "0x1108000432000200142A040200142A040000400A0542006222042200240010400100000000000085",
		INITVAL_05 => "0x1320000001100AA0400A1460205409034020422800238040820A60004400144AA040220108811088",
		INITVAL_06 => "0x06020000121500A044020408810481100A0032130000000280014AA044081042114083004280A410",
		INITVAL_07 => "0x044120422904402042290400100000000AA154AA154AA0440210082004011542214020024081460A",
		INITVAL_08 => "0x100020208000002064120041205000010090A412024090A41204221100950420012A220A4500A421",
		INITVAL_09 => "0x04052142810440A01400044080302A01400004220000214028100A20440204002040020400004400",
		INITVAL_0a => "0x144201140A0042A146A204088110881108010008104500100204400042220A0100048A0000000400",
		INITVAL_0b => "0x0200202402000AA154A20408810012114020B0130402004000044000000510400040030040015420",
		INITVAL_0c => "0x0442800452002300400206232006810740A1542006420110881002004081004A200000020080A402",
		INITVAL_0d => "0x040080A621040010002200600014AA144800102001000144201100804020040A50640802602002A0",
		INITVAL_0e => "0x0120A1442001088014210400213010020AA14028000280040800413120A20029203201040881102A",
		INITVAL_0f => "0x11052050AA154AA1542804008100000000000099132050403300600012001329202E000529202402",
		INITVAL_10 => "0x0049904225040000000012009124090B22104000100010720000413140A0002980041A05012040A1",
		INITVAL_11 => "0x00021000900000900099132100129A0263700099042021429A0242A0000012009132910009904A70",
		INITVAL_12 => "0x1462A152A20A002000030000A024020200A000001200913221142AA0402004032024250008100000",
		INITVAL_13 => "0x0000210621000001002110A210522100080034AA154220000001090020221040811088110880000A",
		INITVAL_14 => "0x1549A044081108804003000001200913203060250000000099006020A0001000302003120320B200",
		INITVAL_15 => "0x14428040881100A040A0114A004A08104520420200085004091008101281144880A6211040003432",
		INITVAL_16 => "0x154AA154A204088104001542A010020208804A200300200280142990B09505295042081040A020AA",
		INITVAL_17 => "0x104020062000410024520A412070020040014A20004820A458064221400004229144A504010050AA",
		INITVAL_18 => "0x120080B0000263904A9810A801041A000350463504630062A20422900202040A0066200242004A21",
		INITVAL_19 => "0x01088110881102000A2006A220140000000120991241307288026380045307012122880105000419",
		INITVAL_1a => "0x01200000981329A0000001209132A30045307225102201141206022014AA15420000AA0B45804232",
		INITVAL_1b => "0x100800028506029010850640200A00110250607900200014AA154AA154901140A04408110AA154A0",
		INITVAL_1c => "0x0122000608040A0052851008000200070A900013000900A0090020A00029102A0010890145900012",
		INITVAL_1d => "0x010201001A014AA15208140A20408814A00150901442011088110881008210085140A000088002A2",
		INITVAL_1e => "0x02083020A00149010A0811252140020520110020002A81000A000850000000400040191000A03005",
		INITVAL_1f => "0x0000901299042331305804AA0004880200A0540A044081108810082000A511013100A0004900300A",
		INITVAL_20 => "0x020080A6390020104A98002800402214000004100340A154901140A0440810400014981002514000",
		INITVAL_21 => "0x13400132A0000000129913492024A90B022044A202492034220B25800422010211005A0248500280",
		INITVAL_22 => "0x00402000000020106010000000A0000A010000030000200000020320108811008140050540014009",
		INITVAL_23 => "0x0000000000000000000000A3200C020E0670E4700CC27000060AC6604C6600C33004720E4660C400"
	)
	port map (
		DIA0 => dmem_write_out(28), DIA1 => dmem_write_out(29),
		DIA2 => dmem_write_out(30), DIA3 => dmem_write_out(31),
		DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
		DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0',
		DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
		DIA16 => '0', DIA17 => '0', 
		DOA0 => dmem_data_read(28), DOA1 => dmem_data_read(29),
		DOA2 => dmem_data_read(30), DOA3 => dmem_data_read(31),
		DOA4 => open, DOA5 => open, DOA6 => open, DOA7 => open,
		DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
		DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
		DOA16 => open, DOA17 => open, 
		ADA0 => '0', ADA1 => '0',
		ADA2 => dmem_addr(2), ADA3 => dmem_addr(3),
		ADA4 => dmem_addr(4), ADA5 => dmem_addr(5),
		ADA6 => dmem_addr(6), ADA7 => dmem_addr(7),
		ADA8 => dmem_addr(8), ADA9 => dmem_addr(9),
		ADA10 => dmem_addr(10), ADA11 => dmem_addr(11),
		ADA12 => dmem_addr(12), ADA13 => dmem_addr(13),
		CEA => dmem_bram_cs, CLKA => not clk, WEA => dmem_write,
		CSA0 => not dmem_byte_sel(3), CSA1 => '0', CSA2 => '0',
		RSTA => '0',

		DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0', 
		DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0', 
		DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
		DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0', 
		DIB16 => '0', DIB17 => '0',
		DOB0 => imem_data_out(28), DOB1 => imem_data_out(29),
		DOB2 => imem_data_out(30), DOB3 => imem_data_out(31),
		DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
		DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
		DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
		DOB16 => open, DOB17 => open, 
		ADB0 => '0', ADB1 => '0',
		ADB2 => imem_addr(2), ADB3 => imem_addr(3),
		ADB4 => imem_addr(4), ADB5 => imem_addr(5),
		ADB6 => imem_addr(6), ADB7 => imem_addr(7),
		ADB8 => imem_addr(8), ADB9 => imem_addr(9),
		ADB10 => imem_addr(10), ADB11 => imem_addr(11),
		ADB12 => imem_addr(12), ADB13 => imem_addr(13),
		CEB => '1', CLKB => not clk, WEB => '0', 
		CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);
	end generate; -- 16k

end Behavioral;
