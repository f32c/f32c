--
-- Copyright 2010 University of Zagreb, Croatia.
--
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions
-- are met:
-- 1. Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimer.
-- 2. Redistributions in binary form must reproduce the above copyright
--    notice, this list of conditions and the following disclaimer in the
--    documentation and/or other materials provided with the distribution.
--
-- THIS SOFTWARE IS PROVIDED BY AUTHOR AND CONTRIBUTORS ``AS IS'' AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
-- IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
-- ARE DISCLAIMED.  IN NO EVENT SHALL AUTHOR OR CONTRIBUTORS BE LIABLE
-- FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL
-- DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS
-- OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
-- HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
-- LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY
-- OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF
-- SUCH DAMAGE.
--

-- $Id: serial.vhd 116 2011-03-28 12:43:12Z marko $

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library xp2;
use xp2.components.all;

entity serial_debug is
	generic (
		clk_divisor: std_logic_vector(15 downto 0)
			-- := x"1458" -- 9600 bps
			:= x"0a2c" -- 19200 bps
			-- := x"0516" -- 38400 bps
			-- := x"0364" -- 57600 bps
			-- := x"01b2" -- 115200 bps
			-- := x"00d9" -- 230400 bps
	);
	port (
		clk: in std_logic;
		rs232_txd: out std_logic;
		trace_addr: out std_logic_vector(5 downto 0);
		trace_data: in std_logic_vector(31 downto 0)
	);
end serial_debug;

architecture Behavioral of serial_debug is
	signal rs232_tick_cnt: std_logic_vector(15 downto 0);
	signal txd: std_logic;
	signal txbitcnt: std_logic_vector(3 downto 0);
	signal txchar, nextchar: std_logic_vector(7 downto 0);
	signal char_tx_done: boolean;
	signal trace_phase: std_logic_vector(3 downto 0);
	signal trace_word: std_logic_vector(31 downto 0);
	signal trace_addr_next: std_logic_vector(5 downto 0);
	signal bram_out: std_logic_vector(7 downto 0);
	signal bram_addr: std_logic_vector(10 downto 0);

begin

	rs232_txd <= txd;
	trace_addr <= trace_addr_next;
	
	debug_rom: DP16KB
	generic map (
	    INITVAL_3F=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
	    INITVAL_3E=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
	    INITVAL_3D=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_3C=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_3B=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_3A=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_39=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_38=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_37=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_36=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_35=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_34=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_33=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_32=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_31=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_30=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2F=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2E=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2D=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2C=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2B=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_2A=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_29=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_28=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_27=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_26=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_25=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_24=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_23=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_22=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_21=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_20=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1F=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1E=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1D=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1C=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1B=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_1A=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_19=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_18=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_17=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_16=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_15=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_14=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_13=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_12=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_11=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_10=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0F=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0E=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0D=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0C=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0B=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_0A=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_09=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_08=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_07=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_06=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_05=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_04=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_03=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_02=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_01=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
            INITVAL_00=> "0x06431060200643106020064310602006431060200643106020064310602006431060200643106020", 
	    -- CSDECODE_B => "111", CSDECODE_A => "000",
	    WRITEMODE_B => "NORMAL", WRITEMODE_A => "NORMAL",
	    GSR => "DISABLED", RESETMODE => "SYNC", 
	    REGMODE_B => "NOREG", REGMODE_A => "NOREG",
	    DATA_WIDTH_B => 9, DATA_WIDTH_A=> 9
	)
	port map (
	    DIA0 => '0', DIA1 => '0', DIA2 => '0', DIA3 => '0',
	    DIA4 => '0', DIA5 => '0', DIA6 => '0', DIA7 => '0',
	    DIA8 => '0', DIA9 => '0', DIA10 => '0', DIA11 => '0', 
	    DIA12 => '0', DIA13 => '0', DIA14 => '0', DIA15 => '0',
	    DIA16 => '0', DIA17 => '0', 
	    DOA0 => bram_out(0), DOA1 => bram_out(1), DOA2 => bram_out(2), DOA3 => bram_out(3),
	    DOA4 => bram_out(4), DOA5 => bram_out(5), DOA6 => bram_out(6), DOA7 => bram_out(7),
	    DOA8 => open, DOA9 => open, DOA10 => open, DOA11 => open,
	    DOA12 => open, DOA13 => open, DOA14 => open, DOA15 => open,
	    DOA16 => open, DOA17 => open, 
	    ADA0 => '0', ADA1 => '0', ADA2 => '0', ADA3 => bram_addr(0),
	    ADA4 => bram_addr(1), ADA5 => bram_addr(2), ADA6 => bram_addr(3), ADA7 => bram_addr(4),
	    ADA8 => bram_addr(5), ADA9 => bram_addr(6), ADA10 => bram_addr(7), ADA11 => bram_addr(8), 
	    ADA12 => bram_addr(9), ADA13 => bram_addr(10),
	    CEA => '1', CLKA => clk, WEA => '0',
	    CSA0 => '0', CSA1 => '0', CSA2 => '0', RSTA => '0', 

	    DIB0 => '0', DIB1 => '0', DIB2 => '0', DIB3 => '0',
	    DIB4 => '0', DIB5 => '0', DIB6 => '0', DIB7 => '0',
	    DIB8 => '0', DIB9 => '0', DIB10 => '0', DIB11 => '0', 
	    DIB12 => '0', DIB13 => '0', DIB14 => '0', DIB15 => '0',
	    DIB16 => '0', DIB17 => '0', 
	    DOB0 => open, DOB1 => open, DOB2 => open, DOB3 => open,
	    DOB4 => open, DOB5 => open, DOB6 => open, DOB7 => open,
	    DOB8 => open, DOB9 => open, DOB10 => open, DOB11 => open,
	    DOB12 => open, DOB13 => open, DOB14 => open, DOB15 => open,
	    DOB16 => open, DOB17 => open,
	    ADB0 => '0', ADB1 => '0', ADB2 => '0', ADB3 => '0',
	    ADB4 => '0', ADB5 => '0', ADB6 => '0', ADB7 => '0',
	    ADB8 => '0', ADB9 => '0', ADB10 => '0', ADB11 => '0', 
	    ADB12 => '0', ADB13 => '0',
	    CEB => '0', CLKB => '0', WEB => '0',
	    CSB0 => '0', CSB1 => '0', CSB2 => '0', RSTB => '0'
	);

	process(clk)
	begin
		if rising_edge(clk) then
		
			-- TX a char, bit by bit
			char_tx_done <= false;
			rs232_tick_cnt <= rs232_tick_cnt - 1;
			if rs232_tick_cnt = "0000" then
				rs232_tick_cnt <= clk_divisor;
				txbitcnt <= txbitcnt + 1;
				txd <= txchar(0);
				txchar <= '1' & txchar(7 downto 1);
				if txbitcnt = "1010" then
					txbitcnt <= "0000";
					txd <= '0'; -- start bit
					txchar <= nextchar;
					char_tx_done <= true;
				end if;
			end if;
			
			-- Fetch new char
			if char_tx_done then
				if trace_phase /= "0000" then
					-- print out trace word in hex one nibble at a time
					trace_phase <= trace_phase - 1;
					if trace_word(31 downto 28) < "1010" then
						nextchar <= "00110000" + trace_word(31 downto 28);
					else
						nextchar <= "01010111" + trace_word(31 downto 28);
					end if;
					trace_word(31 downto 4) <= trace_word(27 downto 0);
				else
					bram_addr <= bram_addr + 1;
					if bram_out(7 downto 6) = "10" then
						-- set new trace addr
						trace_addr_next <= bram_out(5 downto 0);
						nextchar <= x"00";
					elsif bram_out(7 downto 5) = "110" then
						-- fetch new trace word and start printing it out
						trace_word <= trace_data;
						trace_phase <= "1000";
						nextchar <= x"00";
					elsif bram_out(7 downto 5) = "111" then
						-- goto bram address 0
						bram_addr <= "00000000000";
						nextchar <= x"00";
					else
						-- ordinary ASCII character - print it out
						nextchar <= bram_out;
					end if;
				end if;
			end if;
		end if;
	end process;

end Behavioral;
